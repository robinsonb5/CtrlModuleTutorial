-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb9",
     9 => x"d0080b0b",
    10 => x"0bb9d408",
    11 => x"0b0b0bb9",
    12 => x"d8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b9d80c0b",
    16 => x"0b0bb9d4",
    17 => x"0c0b0b0b",
    18 => x"b9d00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb2b0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b9d07080",
    57 => x"c48c278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"51888804",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb9e00c",
    65 => x"9f0bb9e4",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b9e408ff",
    69 => x"05b9e40c",
    70 => x"b9e40880",
    71 => x"25eb38b9",
    72 => x"e008ff05",
    73 => x"b9e00cb9",
    74 => x"e0088025",
    75 => x"d738800b",
    76 => x"b9e40c80",
    77 => x"0bb9e00c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb9e008",
    97 => x"258f3882",
    98 => x"bd2db9e0",
    99 => x"08ff05b9",
   100 => x"e00c82ff",
   101 => x"04b9e008",
   102 => x"b9e40853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b9e008a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b9e4",
   111 => x"088105b9",
   112 => x"e40cb9e4",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb9e40c",
   116 => x"b9e00881",
   117 => x"05b9e00c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b9",
   122 => x"e4088105",
   123 => x"b9e40cb9",
   124 => x"e408a02e",
   125 => x"0981068e",
   126 => x"38800bb9",
   127 => x"e40cb9e0",
   128 => x"088105b9",
   129 => x"e00c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb9e8",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb9e80c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b9",
   169 => x"e8088407",
   170 => x"b9e80c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb5f4",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfecc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b9e80852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b9d00c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"8dc72d80",
   203 => x"518cfa2d",
   204 => x"8cfa2d8c",
   205 => x"fa2d8cfa",
   206 => x"2d70f00c",
   207 => x"70f40c70",
   208 => x"f80c8111",
   209 => x"51907125",
   210 => x"e4388db4",
   211 => x"2d028405",
   212 => x"0d0402fc",
   213 => x"050dec51",
   214 => x"83710c82",
   215 => x"710c0284",
   216 => x"050d0402",
   217 => x"dc050d80",
   218 => x"59810bec",
   219 => x"0c840bec",
   220 => x"0c7a52b9",
   221 => x"ec51a9d3",
   222 => x"2db9d008",
   223 => x"792e80f9",
   224 => x"38b9f008",
   225 => x"79ff1256",
   226 => x"59567379",
   227 => x"2e8b3881",
   228 => x"1874812a",
   229 => x"555873f7",
   230 => x"38f71858",
   231 => x"81598076",
   232 => x"2580d038",
   233 => x"77527351",
   234 => x"848b2dba",
   235 => x"c452b9ec",
   236 => x"51ac922d",
   237 => x"b9d00880",
   238 => x"2e9a38ba",
   239 => x"c45783fc",
   240 => x"55767084",
   241 => x"055808e8",
   242 => x"0cfc1555",
   243 => x"748025f1",
   244 => x"3887db04",
   245 => x"b9d00859",
   246 => x"848056b9",
   247 => x"ec51abe4",
   248 => x"2dfc8016",
   249 => x"81155556",
   250 => x"758024ff",
   251 => x"b7387880",
   252 => x"2e8738b5",
   253 => x"f85187fc",
   254 => x"04b7a451",
   255 => x"8fc32d78",
   256 => x"b9d00c02",
   257 => x"a4050d04",
   258 => x"02f4050d",
   259 => x"810bec0c",
   260 => x"8d952d89",
   261 => x"e42d81f8",
   262 => x"2d83528c",
   263 => x"fa2d8151",
   264 => x"84f02dff",
   265 => x"12527180",
   266 => x"25f13884",
   267 => x"52880bb6",
   268 => x"f00b81b7",
   269 => x"2d880bb6",
   270 => x"fc0b81b7",
   271 => x"2d880bb7",
   272 => x"880b81b7",
   273 => x"2d71ec0c",
   274 => x"b3f85185",
   275 => x"fe2d9cc5",
   276 => x"2da0ec2d",
   277 => x"b9d00880",
   278 => x"2e8638fe",
   279 => x"5288e804",
   280 => x"ff125271",
   281 => x"8024e738",
   282 => x"71802e80",
   283 => x"dc38b490",
   284 => x"5185fe2d",
   285 => x"b4a85186",
   286 => x"e32d86e3",
   287 => x"51b2a72d",
   288 => x"8db42d89",
   289 => x"f02d8fd3",
   290 => x"2db68c0b",
   291 => x"80f52dba",
   292 => x"a4088106",
   293 => x"53537180",
   294 => x"2e853872",
   295 => x"84075372",
   296 => x"fc0cb6f0",
   297 => x"0b80f52d",
   298 => x"f00cb6fc",
   299 => x"0b80f52d",
   300 => x"f40cb788",
   301 => x"0b80f52d",
   302 => x"f80c8652",
   303 => x"b9d00883",
   304 => x"38845271",
   305 => x"ec0c8983",
   306 => x"04b4b451",
   307 => x"85fe2d80",
   308 => x"0bb9d00c",
   309 => x"028c050d",
   310 => x"0471980c",
   311 => x"04ffb008",
   312 => x"b9d00c04",
   313 => x"810bffb0",
   314 => x"0c04800b",
   315 => x"ffb00c04",
   316 => x"02f4050d",
   317 => x"8af204b9",
   318 => x"d00881f0",
   319 => x"2e098106",
   320 => x"8938810b",
   321 => x"b8880c8a",
   322 => x"f204b9d0",
   323 => x"0881e02e",
   324 => x"09810689",
   325 => x"38810bb8",
   326 => x"8c0c8af2",
   327 => x"04b9d008",
   328 => x"52b88c08",
   329 => x"802e8838",
   330 => x"b9d00881",
   331 => x"80055271",
   332 => x"842c728f",
   333 => x"065353b8",
   334 => x"8808802e",
   335 => x"99387284",
   336 => x"29b7c805",
   337 => x"72138171",
   338 => x"2b700973",
   339 => x"0806730c",
   340 => x"5153538a",
   341 => x"e8047284",
   342 => x"29b7c805",
   343 => x"72138371",
   344 => x"2b720807",
   345 => x"720c5353",
   346 => x"800bb88c",
   347 => x"0c800bb8",
   348 => x"880cb9f8",
   349 => x"518bf32d",
   350 => x"b9d008ff",
   351 => x"24fef838",
   352 => x"800bb9d0",
   353 => x"0c028c05",
   354 => x"0d0402f8",
   355 => x"050db7c8",
   356 => x"528f5180",
   357 => x"72708405",
   358 => x"540cff11",
   359 => x"51708025",
   360 => x"f2380288",
   361 => x"050d0402",
   362 => x"f0050d75",
   363 => x"5189ea2d",
   364 => x"70822cfc",
   365 => x"06b7c811",
   366 => x"72109e06",
   367 => x"71087072",
   368 => x"2a708306",
   369 => x"82742b70",
   370 => x"09740676",
   371 => x"0c545156",
   372 => x"57535153",
   373 => x"89e42d71",
   374 => x"b9d00c02",
   375 => x"90050d04",
   376 => x"02fc050d",
   377 => x"72518071",
   378 => x"0c800b84",
   379 => x"120c0284",
   380 => x"050d0402",
   381 => x"f0050d75",
   382 => x"70088412",
   383 => x"08535353",
   384 => x"ff547171",
   385 => x"2ea83889",
   386 => x"ea2d8413",
   387 => x"08708429",
   388 => x"14881170",
   389 => x"087081ff",
   390 => x"06841808",
   391 => x"81118706",
   392 => x"841a0c53",
   393 => x"51555151",
   394 => x"5189e42d",
   395 => x"715473b9",
   396 => x"d00c0290",
   397 => x"050d0402",
   398 => x"f8050d89",
   399 => x"ea2de008",
   400 => x"708b2a70",
   401 => x"81065152",
   402 => x"5270802e",
   403 => x"9d38b9f8",
   404 => x"08708429",
   405 => x"ba800573",
   406 => x"81ff0671",
   407 => x"0c5151b9",
   408 => x"f8088111",
   409 => x"8706b9f8",
   410 => x"0c51800b",
   411 => x"baa00c89",
   412 => x"dd2d89e4",
   413 => x"2d028805",
   414 => x"0d0402fc",
   415 => x"050d89ea",
   416 => x"2d810bba",
   417 => x"a00c89e4",
   418 => x"2dbaa008",
   419 => x"5170fa38",
   420 => x"0284050d",
   421 => x"0402fc05",
   422 => x"0db9f851",
   423 => x"8be02d8b",
   424 => x"8a2d8cb7",
   425 => x"5189d92d",
   426 => x"0284050d",
   427 => x"04bab008",
   428 => x"b9d00c04",
   429 => x"02fc050d",
   430 => x"810bb890",
   431 => x"0c815184",
   432 => x"f02d0284",
   433 => x"050d0402",
   434 => x"fc050d8d",
   435 => x"d10489f0",
   436 => x"2d87518b",
   437 => x"a72db9d0",
   438 => x"08f43880",
   439 => x"da518ba7",
   440 => x"2db9d008",
   441 => x"e938b9d0",
   442 => x"08b8900c",
   443 => x"b9d00851",
   444 => x"84f02d02",
   445 => x"84050d04",
   446 => x"02ec050d",
   447 => x"76548052",
   448 => x"870b8815",
   449 => x"80f52d56",
   450 => x"53747224",
   451 => x"8338a053",
   452 => x"725182f9",
   453 => x"2d81128b",
   454 => x"1580f52d",
   455 => x"54527272",
   456 => x"25de3802",
   457 => x"94050d04",
   458 => x"02f0050d",
   459 => x"bab00854",
   460 => x"81f82d80",
   461 => x"0bbab40c",
   462 => x"7308802e",
   463 => x"81803882",
   464 => x"0bb9e40c",
   465 => x"bab4088f",
   466 => x"06b9e00c",
   467 => x"73085271",
   468 => x"832e9638",
   469 => x"71832689",
   470 => x"3871812e",
   471 => x"af388fa9",
   472 => x"0471852e",
   473 => x"9f388fa9",
   474 => x"04881480",
   475 => x"f52d8415",
   476 => x"08b4c853",
   477 => x"545285fe",
   478 => x"2d718429",
   479 => x"13700852",
   480 => x"528fad04",
   481 => x"73518df8",
   482 => x"2d8fa904",
   483 => x"baa40888",
   484 => x"15082c70",
   485 => x"81065152",
   486 => x"71802e87",
   487 => x"38b4cc51",
   488 => x"8fa604b4",
   489 => x"d05185fe",
   490 => x"2d841408",
   491 => x"5185fe2d",
   492 => x"bab40881",
   493 => x"05bab40c",
   494 => x"8c14548e",
   495 => x"b8040290",
   496 => x"050d0471",
   497 => x"bab00c8e",
   498 => x"a82dbab4",
   499 => x"08ff05ba",
   500 => x"b80c0402",
   501 => x"e8050dba",
   502 => x"b008babc",
   503 => x"08575587",
   504 => x"518ba72d",
   505 => x"b9d00881",
   506 => x"2a708106",
   507 => x"51527180",
   508 => x"2ea0388f",
   509 => x"f90489f0",
   510 => x"2d87518b",
   511 => x"a72db9d0",
   512 => x"08f438b8",
   513 => x"90088132",
   514 => x"70b8900c",
   515 => x"70525284",
   516 => x"f02d800b",
   517 => x"baa80c80",
   518 => x"0bbaac0c",
   519 => x"b8900882",
   520 => x"dd3880da",
   521 => x"518ba72d",
   522 => x"b9d00880",
   523 => x"2e8a38ba",
   524 => x"a8088180",
   525 => x"07baa80c",
   526 => x"80d9518b",
   527 => x"a72db9d0",
   528 => x"08802e8a",
   529 => x"38baa808",
   530 => x"80c007ba",
   531 => x"a80c8194",
   532 => x"518ba72d",
   533 => x"b9d00880",
   534 => x"2e8938ba",
   535 => x"a8089007",
   536 => x"baa80c81",
   537 => x"91518ba7",
   538 => x"2db9d008",
   539 => x"802e8938",
   540 => x"baa808a0",
   541 => x"07baa80c",
   542 => x"81f5518b",
   543 => x"a72db9d0",
   544 => x"08802e89",
   545 => x"38baa808",
   546 => x"8107baa8",
   547 => x"0c81f251",
   548 => x"8ba72db9",
   549 => x"d008802e",
   550 => x"8938baa8",
   551 => x"088207ba",
   552 => x"a80c81eb",
   553 => x"518ba72d",
   554 => x"b9d00880",
   555 => x"2e8938ba",
   556 => x"a8088407",
   557 => x"baa80c81",
   558 => x"f4518ba7",
   559 => x"2db9d008",
   560 => x"802e8938",
   561 => x"baa80888",
   562 => x"07baa80c",
   563 => x"80d8518b",
   564 => x"a72db9d0",
   565 => x"08802e8a",
   566 => x"38baac08",
   567 => x"818007ba",
   568 => x"ac0c9251",
   569 => x"8ba72db9",
   570 => x"d008802e",
   571 => x"8a38baac",
   572 => x"0880c007",
   573 => x"baac0c94",
   574 => x"518ba72d",
   575 => x"b9d00880",
   576 => x"2e8938ba",
   577 => x"ac089007",
   578 => x"baac0c91",
   579 => x"518ba72d",
   580 => x"b9d00880",
   581 => x"2e8938ba",
   582 => x"ac08a007",
   583 => x"baac0c9d",
   584 => x"518ba72d",
   585 => x"b9d00880",
   586 => x"2e8938ba",
   587 => x"ac088107",
   588 => x"baac0c9b",
   589 => x"518ba72d",
   590 => x"b9d00880",
   591 => x"2e8938ba",
   592 => x"ac088207",
   593 => x"baac0c9c",
   594 => x"518ba72d",
   595 => x"b9d00880",
   596 => x"2e8938ba",
   597 => x"ac088407",
   598 => x"baac0ca3",
   599 => x"518ba72d",
   600 => x"b9d00880",
   601 => x"2e8938ba",
   602 => x"ac088807",
   603 => x"baac0c81",
   604 => x"fd518ba7",
   605 => x"2d81fa51",
   606 => x"8ba72d98",
   607 => x"af0481f5",
   608 => x"518ba72d",
   609 => x"b9d00881",
   610 => x"2a708106",
   611 => x"51527180",
   612 => x"2eaf38ba",
   613 => x"b8085271",
   614 => x"802e8938",
   615 => x"ff12bab8",
   616 => x"0c93c104",
   617 => x"bab40810",
   618 => x"bab40805",
   619 => x"70842916",
   620 => x"51528812",
   621 => x"08802e89",
   622 => x"38ff5188",
   623 => x"12085271",
   624 => x"2d81f251",
   625 => x"8ba72db9",
   626 => x"d008812a",
   627 => x"70810651",
   628 => x"5271802e",
   629 => x"b138bab4",
   630 => x"08ff11ba",
   631 => x"b8085653",
   632 => x"53737225",
   633 => x"89388114",
   634 => x"bab80c94",
   635 => x"86047210",
   636 => x"13708429",
   637 => x"16515288",
   638 => x"1208802e",
   639 => x"8938fe51",
   640 => x"88120852",
   641 => x"712d81fd",
   642 => x"518ba72d",
   643 => x"b9d00881",
   644 => x"2a708106",
   645 => x"51527180",
   646 => x"2ead38ba",
   647 => x"b808802e",
   648 => x"8938800b",
   649 => x"bab80c94",
   650 => x"c704bab4",
   651 => x"0810bab4",
   652 => x"08057084",
   653 => x"29165152",
   654 => x"88120880",
   655 => x"2e8938fd",
   656 => x"51881208",
   657 => x"52712d81",
   658 => x"fa518ba7",
   659 => x"2db9d008",
   660 => x"812a7081",
   661 => x"06515271",
   662 => x"802eae38",
   663 => x"bab408ff",
   664 => x"115452ba",
   665 => x"b8087325",
   666 => x"883872ba",
   667 => x"b80c9589",
   668 => x"04711012",
   669 => x"70842916",
   670 => x"51528812",
   671 => x"08802e89",
   672 => x"38fc5188",
   673 => x"12085271",
   674 => x"2dbab808",
   675 => x"70535473",
   676 => x"802e8a38",
   677 => x"8c15ff15",
   678 => x"5555958f",
   679 => x"04820bb9",
   680 => x"e40c718f",
   681 => x"06b9e00c",
   682 => x"81eb518b",
   683 => x"a72db9d0",
   684 => x"08812a70",
   685 => x"81065152",
   686 => x"71802ead",
   687 => x"38740885",
   688 => x"2e098106",
   689 => x"a4388815",
   690 => x"80f52dff",
   691 => x"05527188",
   692 => x"1681b72d",
   693 => x"71982b52",
   694 => x"71802588",
   695 => x"38800b88",
   696 => x"1681b72d",
   697 => x"74518df8",
   698 => x"2d81f451",
   699 => x"8ba72db9",
   700 => x"d008812a",
   701 => x"70810651",
   702 => x"5271802e",
   703 => x"b3387408",
   704 => x"852e0981",
   705 => x"06aa3888",
   706 => x"1580f52d",
   707 => x"81055271",
   708 => x"881681b7",
   709 => x"2d7181ff",
   710 => x"068b1680",
   711 => x"f52d5452",
   712 => x"72722787",
   713 => x"38728816",
   714 => x"81b72d74",
   715 => x"518df82d",
   716 => x"80da518b",
   717 => x"a72db9d0",
   718 => x"08812a70",
   719 => x"81065152",
   720 => x"71802e81",
   721 => x"a638bab0",
   722 => x"08bab808",
   723 => x"55537380",
   724 => x"2e8a388c",
   725 => x"13ff1555",
   726 => x"5396ce04",
   727 => x"72085271",
   728 => x"822ea638",
   729 => x"71822689",
   730 => x"3871812e",
   731 => x"a93897eb",
   732 => x"0471832e",
   733 => x"b1387184",
   734 => x"2e098106",
   735 => x"80ed3888",
   736 => x"1308518f",
   737 => x"c32d97eb",
   738 => x"04bab808",
   739 => x"51881308",
   740 => x"52712d97",
   741 => x"eb04810b",
   742 => x"8814082b",
   743 => x"baa40832",
   744 => x"baa40c97",
   745 => x"c1048813",
   746 => x"80f52d81",
   747 => x"058b1480",
   748 => x"f52d5354",
   749 => x"71742483",
   750 => x"38805473",
   751 => x"881481b7",
   752 => x"2d8ea82d",
   753 => x"97eb0475",
   754 => x"08802ea2",
   755 => x"38750851",
   756 => x"8ba72db9",
   757 => x"d0088106",
   758 => x"5271802e",
   759 => x"8b38bab8",
   760 => x"08518416",
   761 => x"0852712d",
   762 => x"88165675",
   763 => x"da388054",
   764 => x"800bb9e4",
   765 => x"0c738f06",
   766 => x"b9e00ca0",
   767 => x"5273bab8",
   768 => x"082e0981",
   769 => x"069838ba",
   770 => x"b408ff05",
   771 => x"74327009",
   772 => x"81057072",
   773 => x"079f2a91",
   774 => x"71315151",
   775 => x"53537151",
   776 => x"82f92d81",
   777 => x"14548e74",
   778 => x"25c638b8",
   779 => x"90085271",
   780 => x"b9d00c02",
   781 => x"98050d04",
   782 => x"02f4050d",
   783 => x"d45281ff",
   784 => x"720c7108",
   785 => x"5381ff72",
   786 => x"0c72882b",
   787 => x"83fe8006",
   788 => x"72087081",
   789 => x"ff065152",
   790 => x"5381ff72",
   791 => x"0c727107",
   792 => x"882b7208",
   793 => x"7081ff06",
   794 => x"51525381",
   795 => x"ff720c72",
   796 => x"7107882b",
   797 => x"72087081",
   798 => x"ff067207",
   799 => x"b9d00c52",
   800 => x"53028c05",
   801 => x"0d0402f4",
   802 => x"050d7476",
   803 => x"7181ff06",
   804 => x"d40c5353",
   805 => x"bac00885",
   806 => x"3871892b",
   807 => x"5271982a",
   808 => x"d40c7190",
   809 => x"2a7081ff",
   810 => x"06d40c51",
   811 => x"71882a70",
   812 => x"81ff06d4",
   813 => x"0c517181",
   814 => x"ff06d40c",
   815 => x"72902a70",
   816 => x"81ff06d4",
   817 => x"0c51d408",
   818 => x"7081ff06",
   819 => x"515182b8",
   820 => x"bf527081",
   821 => x"ff2e0981",
   822 => x"06943881",
   823 => x"ff0bd40c",
   824 => x"d4087081",
   825 => x"ff06ff14",
   826 => x"54515171",
   827 => x"e53870b9",
   828 => x"d00c028c",
   829 => x"050d0402",
   830 => x"fc050d81",
   831 => x"c75181ff",
   832 => x"0bd40cff",
   833 => x"11517080",
   834 => x"25f43802",
   835 => x"84050d04",
   836 => x"02f0050d",
   837 => x"99f72d8f",
   838 => x"cf538052",
   839 => x"87fc80f7",
   840 => x"5199862d",
   841 => x"b9d00854",
   842 => x"b9d00881",
   843 => x"2e098106",
   844 => x"a33881ff",
   845 => x"0bd40c82",
   846 => x"0a52849c",
   847 => x"80e95199",
   848 => x"862db9d0",
   849 => x"088b3881",
   850 => x"ff0bd40c",
   851 => x"73539ada",
   852 => x"0499f72d",
   853 => x"ff135372",
   854 => x"c13872b9",
   855 => x"d00c0290",
   856 => x"050d0402",
   857 => x"f4050d81",
   858 => x"ff0bd40c",
   859 => x"93538052",
   860 => x"87fc80c1",
   861 => x"5199862d",
   862 => x"b9d0088b",
   863 => x"3881ff0b",
   864 => x"d40c8153",
   865 => x"9b900499",
   866 => x"f72dff13",
   867 => x"5372df38",
   868 => x"72b9d00c",
   869 => x"028c050d",
   870 => x"0402f005",
   871 => x"0d99f72d",
   872 => x"83aa5284",
   873 => x"9c80c851",
   874 => x"99862db9",
   875 => x"d008812e",
   876 => x"09810692",
   877 => x"3898b82d",
   878 => x"b9d00883",
   879 => x"ffff0653",
   880 => x"7283aa2e",
   881 => x"97389ae3",
   882 => x"2d9bd704",
   883 => x"81549cbc",
   884 => x"04b4d451",
   885 => x"85fe2d80",
   886 => x"549cbc04",
   887 => x"81ff0bd4",
   888 => x"0cb1539a",
   889 => x"902db9d0",
   890 => x"08802e80",
   891 => x"c0388052",
   892 => x"87fc80fa",
   893 => x"5199862d",
   894 => x"b9d008b1",
   895 => x"3881ff0b",
   896 => x"d40cd408",
   897 => x"5381ff0b",
   898 => x"d40c81ff",
   899 => x"0bd40c81",
   900 => x"ff0bd40c",
   901 => x"81ff0bd4",
   902 => x"0c72862a",
   903 => x"708106b9",
   904 => x"d0085651",
   905 => x"5372802e",
   906 => x"93389bcc",
   907 => x"0472822e",
   908 => x"ff9f38ff",
   909 => x"135372ff",
   910 => x"aa387254",
   911 => x"73b9d00c",
   912 => x"0290050d",
   913 => x"0402f005",
   914 => x"0d810bba",
   915 => x"c00c8454",
   916 => x"d008708f",
   917 => x"2a708106",
   918 => x"51515372",
   919 => x"f33872d0",
   920 => x"0c99f72d",
   921 => x"b4e45185",
   922 => x"fe2dd008",
   923 => x"708f2a70",
   924 => x"81065151",
   925 => x"5372f338",
   926 => x"810bd00c",
   927 => x"b1538052",
   928 => x"84d480c0",
   929 => x"5199862d",
   930 => x"b9d00881",
   931 => x"2ea13872",
   932 => x"822e0981",
   933 => x"068c38b4",
   934 => x"f05185fe",
   935 => x"2d80539d",
   936 => x"e404ff13",
   937 => x"5372d738",
   938 => x"ff145473",
   939 => x"ffa2389b",
   940 => x"992db9d0",
   941 => x"08bac00c",
   942 => x"b9d0088b",
   943 => x"38815287",
   944 => x"fc80d051",
   945 => x"99862d81",
   946 => x"ff0bd40c",
   947 => x"d008708f",
   948 => x"2a708106",
   949 => x"51515372",
   950 => x"f33872d0",
   951 => x"0c81ff0b",
   952 => x"d40c8153",
   953 => x"72b9d00c",
   954 => x"0290050d",
   955 => x"0402e805",
   956 => x"0d785580",
   957 => x"5681ff0b",
   958 => x"d40cd008",
   959 => x"708f2a70",
   960 => x"81065151",
   961 => x"5372f338",
   962 => x"82810bd0",
   963 => x"0c81ff0b",
   964 => x"d40c7752",
   965 => x"87fc80d1",
   966 => x"5199862d",
   967 => x"80dbc6df",
   968 => x"54b9d008",
   969 => x"802e8a38",
   970 => x"b5985185",
   971 => x"fe2d9f84",
   972 => x"0481ff0b",
   973 => x"d40cd408",
   974 => x"7081ff06",
   975 => x"51537281",
   976 => x"fe2e0981",
   977 => x"069d3880",
   978 => x"ff5398b8",
   979 => x"2db9d008",
   980 => x"75708405",
   981 => x"570cff13",
   982 => x"53728025",
   983 => x"ed388156",
   984 => x"9ee904ff",
   985 => x"145473c9",
   986 => x"3881ff0b",
   987 => x"d40c81ff",
   988 => x"0bd40cd0",
   989 => x"08708f2a",
   990 => x"70810651",
   991 => x"515372f3",
   992 => x"3872d00c",
   993 => x"75b9d00c",
   994 => x"0298050d",
   995 => x"0402e805",
   996 => x"0d77797b",
   997 => x"58555580",
   998 => x"53727625",
   999 => x"a3387470",
  1000 => x"81055680",
  1001 => x"f52d7470",
  1002 => x"81055680",
  1003 => x"f52d5252",
  1004 => x"71712e86",
  1005 => x"3881519f",
  1006 => x"c2048113",
  1007 => x"539f9904",
  1008 => x"805170b9",
  1009 => x"d00c0298",
  1010 => x"050d0402",
  1011 => x"ec050d76",
  1012 => x"5574802e",
  1013 => x"be389a15",
  1014 => x"80e02d51",
  1015 => x"aceb2db9",
  1016 => x"d008b9d0",
  1017 => x"0880c0f4",
  1018 => x"0cb9d008",
  1019 => x"545480c0",
  1020 => x"d008802e",
  1021 => x"99389415",
  1022 => x"80e02d51",
  1023 => x"aceb2db9",
  1024 => x"d008902b",
  1025 => x"83fff00a",
  1026 => x"06707507",
  1027 => x"51537280",
  1028 => x"c0f40c80",
  1029 => x"c0f40853",
  1030 => x"72802e9d",
  1031 => x"3880c0c8",
  1032 => x"08fe1471",
  1033 => x"2980c0dc",
  1034 => x"080580c0",
  1035 => x"f80c7084",
  1036 => x"2b80c0d4",
  1037 => x"0c54a0e7",
  1038 => x"0480c0e0",
  1039 => x"0880c0f4",
  1040 => x"0c80c0e4",
  1041 => x"0880c0f8",
  1042 => x"0c80c0d0",
  1043 => x"08802e8b",
  1044 => x"3880c0c8",
  1045 => x"08842b53",
  1046 => x"a0e20480",
  1047 => x"c0e80884",
  1048 => x"2b537280",
  1049 => x"c0d40c02",
  1050 => x"94050d04",
  1051 => x"02d8050d",
  1052 => x"800b80c0",
  1053 => x"d00cbac4",
  1054 => x"5280519d",
  1055 => x"ed2db9d0",
  1056 => x"0854b9d0",
  1057 => x"088c38b5",
  1058 => x"a85185fe",
  1059 => x"2d7355a6",
  1060 => x"a6048056",
  1061 => x"810b80c0",
  1062 => x"fc0c8853",
  1063 => x"b5b452ba",
  1064 => x"fa519f8d",
  1065 => x"2db9d008",
  1066 => x"762e0981",
  1067 => x"068838b9",
  1068 => x"d00880c0",
  1069 => x"fc0c8853",
  1070 => x"b5c052bb",
  1071 => x"96519f8d",
  1072 => x"2db9d008",
  1073 => x"8838b9d0",
  1074 => x"0880c0fc",
  1075 => x"0c80c0fc",
  1076 => x"08802e80",
  1077 => x"f638be8a",
  1078 => x"0b80f52d",
  1079 => x"be8b0b80",
  1080 => x"f52d7198",
  1081 => x"2b71902b",
  1082 => x"07be8c0b",
  1083 => x"80f52d70",
  1084 => x"882b7207",
  1085 => x"be8d0b80",
  1086 => x"f52d7107",
  1087 => x"bec20b80",
  1088 => x"f52dbec3",
  1089 => x"0b80f52d",
  1090 => x"71882b07",
  1091 => x"535f5452",
  1092 => x"5a565755",
  1093 => x"7381abaa",
  1094 => x"2e098106",
  1095 => x"8d387551",
  1096 => x"acbb2db9",
  1097 => x"d00856a2",
  1098 => x"b7047382",
  1099 => x"d4d52e87",
  1100 => x"38b5cc51",
  1101 => x"a2f904ba",
  1102 => x"c4527551",
  1103 => x"9ded2db9",
  1104 => x"d00855b9",
  1105 => x"d008802e",
  1106 => x"83dc3888",
  1107 => x"53b5c052",
  1108 => x"bb96519f",
  1109 => x"8d2db9d0",
  1110 => x"088a3881",
  1111 => x"0b80c0d0",
  1112 => x"0ca2ff04",
  1113 => x"8853b5b4",
  1114 => x"52bafa51",
  1115 => x"9f8d2db9",
  1116 => x"d008802e",
  1117 => x"8a38b5e0",
  1118 => x"5185fe2d",
  1119 => x"a3d904be",
  1120 => x"c20b80f5",
  1121 => x"2d547380",
  1122 => x"d52e0981",
  1123 => x"0680ca38",
  1124 => x"bec30b80",
  1125 => x"f52d5473",
  1126 => x"81aa2e09",
  1127 => x"8106ba38",
  1128 => x"800bbac4",
  1129 => x"0b80f52d",
  1130 => x"56547481",
  1131 => x"e92e8338",
  1132 => x"81547481",
  1133 => x"eb2e8c38",
  1134 => x"80557375",
  1135 => x"2e098106",
  1136 => x"82e438ba",
  1137 => x"cf0b80f5",
  1138 => x"2d55748d",
  1139 => x"38bad00b",
  1140 => x"80f52d54",
  1141 => x"73822e86",
  1142 => x"388055a6",
  1143 => x"a604bad1",
  1144 => x"0b80f52d",
  1145 => x"7080c0c8",
  1146 => x"0cff0580",
  1147 => x"c0cc0cba",
  1148 => x"d20b80f5",
  1149 => x"2dbad30b",
  1150 => x"80f52d58",
  1151 => x"76057782",
  1152 => x"80290570",
  1153 => x"80c0d80c",
  1154 => x"bad40b80",
  1155 => x"f52d7080",
  1156 => x"c0ec0c80",
  1157 => x"c0d00859",
  1158 => x"57587680",
  1159 => x"2e81ac38",
  1160 => x"8853b5c0",
  1161 => x"52bb9651",
  1162 => x"9f8d2db9",
  1163 => x"d00881f6",
  1164 => x"3880c0c8",
  1165 => x"0870842b",
  1166 => x"80c0d40c",
  1167 => x"7080c0e8",
  1168 => x"0cbae90b",
  1169 => x"80f52dba",
  1170 => x"e80b80f5",
  1171 => x"2d718280",
  1172 => x"2905baea",
  1173 => x"0b80f52d",
  1174 => x"70848080",
  1175 => x"2912baeb",
  1176 => x"0b80f52d",
  1177 => x"7081800a",
  1178 => x"29127080",
  1179 => x"c0f00c80",
  1180 => x"c0ec0871",
  1181 => x"2980c0d8",
  1182 => x"08057080",
  1183 => x"c0dc0cba",
  1184 => x"f10b80f5",
  1185 => x"2dbaf00b",
  1186 => x"80f52d71",
  1187 => x"82802905",
  1188 => x"baf20b80",
  1189 => x"f52d7084",
  1190 => x"80802912",
  1191 => x"baf30b80",
  1192 => x"f52d7098",
  1193 => x"2b81f00a",
  1194 => x"06720570",
  1195 => x"80c0e00c",
  1196 => x"fe117e29",
  1197 => x"770580c0",
  1198 => x"e40c5259",
  1199 => x"5243545e",
  1200 => x"51525952",
  1201 => x"5d575957",
  1202 => x"a69f04ba",
  1203 => x"d60b80f5",
  1204 => x"2dbad50b",
  1205 => x"80f52d71",
  1206 => x"82802905",
  1207 => x"7080c0d4",
  1208 => x"0c70a029",
  1209 => x"83ff0570",
  1210 => x"892a7080",
  1211 => x"c0e80cba",
  1212 => x"db0b80f5",
  1213 => x"2dbada0b",
  1214 => x"80f52d71",
  1215 => x"82802905",
  1216 => x"7080c0f0",
  1217 => x"0c7b7129",
  1218 => x"1e7080c0",
  1219 => x"e40c7d80",
  1220 => x"c0e00c73",
  1221 => x"0580c0dc",
  1222 => x"0c555e51",
  1223 => x"51555580",
  1224 => x"519fcb2d",
  1225 => x"815574b9",
  1226 => x"d00c02a8",
  1227 => x"050d0402",
  1228 => x"ec050d76",
  1229 => x"70872c71",
  1230 => x"80ff0655",
  1231 => x"565480c0",
  1232 => x"d0088a38",
  1233 => x"73882c74",
  1234 => x"81ff0654",
  1235 => x"55bac452",
  1236 => x"80c0d808",
  1237 => x"15519ded",
  1238 => x"2db9d008",
  1239 => x"54b9d008",
  1240 => x"802eb438",
  1241 => x"80c0d008",
  1242 => x"802e9838",
  1243 => x"728429ba",
  1244 => x"c4057008",
  1245 => x"5253acbb",
  1246 => x"2db9d008",
  1247 => x"f00a0653",
  1248 => x"a7950472",
  1249 => x"10bac405",
  1250 => x"7080e02d",
  1251 => x"5253aceb",
  1252 => x"2db9d008",
  1253 => x"53725473",
  1254 => x"b9d00c02",
  1255 => x"94050d04",
  1256 => x"02e0050d",
  1257 => x"7970842c",
  1258 => x"80c0f808",
  1259 => x"05718f06",
  1260 => x"52555372",
  1261 => x"8938bac4",
  1262 => x"5273519d",
  1263 => x"ed2d72a0",
  1264 => x"29bac405",
  1265 => x"54807480",
  1266 => x"f52d5653",
  1267 => x"74732e83",
  1268 => x"38815374",
  1269 => x"81e52e81",
  1270 => x"ef388170",
  1271 => x"74065458",
  1272 => x"72802e81",
  1273 => x"e3388b14",
  1274 => x"80f52d70",
  1275 => x"832a7906",
  1276 => x"58567698",
  1277 => x"38b89408",
  1278 => x"53728838",
  1279 => x"72bec40b",
  1280 => x"81b72d76",
  1281 => x"b8940c73",
  1282 => x"53a9ca04",
  1283 => x"758f2e09",
  1284 => x"810681b4",
  1285 => x"38749f06",
  1286 => x"8d29beb7",
  1287 => x"11515381",
  1288 => x"1480f52d",
  1289 => x"73708105",
  1290 => x"5581b72d",
  1291 => x"831480f5",
  1292 => x"2d737081",
  1293 => x"055581b7",
  1294 => x"2d851480",
  1295 => x"f52d7370",
  1296 => x"81055581",
  1297 => x"b72d8714",
  1298 => x"80f52d73",
  1299 => x"70810555",
  1300 => x"81b72d89",
  1301 => x"1480f52d",
  1302 => x"73708105",
  1303 => x"5581b72d",
  1304 => x"8e1480f5",
  1305 => x"2d737081",
  1306 => x"055581b7",
  1307 => x"2d901480",
  1308 => x"f52d7370",
  1309 => x"81055581",
  1310 => x"b72d9214",
  1311 => x"80f52d73",
  1312 => x"70810555",
  1313 => x"81b72d94",
  1314 => x"1480f52d",
  1315 => x"73708105",
  1316 => x"5581b72d",
  1317 => x"961480f5",
  1318 => x"2d737081",
  1319 => x"055581b7",
  1320 => x"2d981480",
  1321 => x"f52d7370",
  1322 => x"81055581",
  1323 => x"b72d9c14",
  1324 => x"80f52d73",
  1325 => x"70810555",
  1326 => x"81b72d9e",
  1327 => x"1480f52d",
  1328 => x"7381b72d",
  1329 => x"77b8940c",
  1330 => x"805372b9",
  1331 => x"d00c02a0",
  1332 => x"050d0402",
  1333 => x"cc050d7e",
  1334 => x"605e5a80",
  1335 => x"0b80c0f4",
  1336 => x"0880c0f8",
  1337 => x"08595c56",
  1338 => x"805880c0",
  1339 => x"d408782e",
  1340 => x"81b03877",
  1341 => x"8f06a017",
  1342 => x"5754738f",
  1343 => x"38bac452",
  1344 => x"76518117",
  1345 => x"579ded2d",
  1346 => x"bac45680",
  1347 => x"7680f52d",
  1348 => x"56547474",
  1349 => x"2e833881",
  1350 => x"547481e5",
  1351 => x"2e80f738",
  1352 => x"81707506",
  1353 => x"555c7380",
  1354 => x"2e80eb38",
  1355 => x"8b1680f5",
  1356 => x"2d980659",
  1357 => x"7880df38",
  1358 => x"8b537c52",
  1359 => x"75519f8d",
  1360 => x"2db9d008",
  1361 => x"80d0389c",
  1362 => x"160851ac",
  1363 => x"bb2db9d0",
  1364 => x"08841b0c",
  1365 => x"9a1680e0",
  1366 => x"2d51aceb",
  1367 => x"2db9d008",
  1368 => x"b9d00888",
  1369 => x"1c0cb9d0",
  1370 => x"08555580",
  1371 => x"c0d00880",
  1372 => x"2e983894",
  1373 => x"1680e02d",
  1374 => x"51aceb2d",
  1375 => x"b9d00890",
  1376 => x"2b83fff0",
  1377 => x"0a067016",
  1378 => x"51547388",
  1379 => x"1b0c787a",
  1380 => x"0c7b54ab",
  1381 => x"db048118",
  1382 => x"5880c0d4",
  1383 => x"087826fe",
  1384 => x"d23880c0",
  1385 => x"d008802e",
  1386 => x"b0387a51",
  1387 => x"a6af2db9",
  1388 => x"d008b9d0",
  1389 => x"0880ffff",
  1390 => x"fff80655",
  1391 => x"5b7380ff",
  1392 => x"fffff82e",
  1393 => x"9438b9d0",
  1394 => x"08fe0580",
  1395 => x"c0c80829",
  1396 => x"80c0dc08",
  1397 => x"0557a9e8",
  1398 => x"04805473",
  1399 => x"b9d00c02",
  1400 => x"b4050d04",
  1401 => x"02f4050d",
  1402 => x"74700881",
  1403 => x"05710c70",
  1404 => x"0880c0cc",
  1405 => x"08065353",
  1406 => x"718e3888",
  1407 => x"130851a6",
  1408 => x"af2db9d0",
  1409 => x"0888140c",
  1410 => x"810bb9d0",
  1411 => x"0c028c05",
  1412 => x"0d0402f0",
  1413 => x"050d7588",
  1414 => x"1108fe05",
  1415 => x"80c0c808",
  1416 => x"2980c0dc",
  1417 => x"08117208",
  1418 => x"80c0cc08",
  1419 => x"06057955",
  1420 => x"5354549d",
  1421 => x"ed2d0290",
  1422 => x"050d0402",
  1423 => x"f4050d74",
  1424 => x"70882a83",
  1425 => x"fe800670",
  1426 => x"72982a07",
  1427 => x"72882b87",
  1428 => x"fc808006",
  1429 => x"73982b81",
  1430 => x"f00a0671",
  1431 => x"730707b9",
  1432 => x"d00c5651",
  1433 => x"5351028c",
  1434 => x"050d0402",
  1435 => x"f8050d02",
  1436 => x"8e0580f5",
  1437 => x"2d74882b",
  1438 => x"077083ff",
  1439 => x"ff06b9d0",
  1440 => x"0c510288",
  1441 => x"050d0402",
  1442 => x"f4050d74",
  1443 => x"76785354",
  1444 => x"52807125",
  1445 => x"97387270",
  1446 => x"81055480",
  1447 => x"f52d7270",
  1448 => x"81055481",
  1449 => x"b72dff11",
  1450 => x"5170eb38",
  1451 => x"807281b7",
  1452 => x"2d028c05",
  1453 => x"0d0402e8",
  1454 => x"050d7756",
  1455 => x"80705654",
  1456 => x"737624b3",
  1457 => x"3880c0d4",
  1458 => x"08742eab",
  1459 => x"387351a7",
  1460 => x"a02db9d0",
  1461 => x"08b9d008",
  1462 => x"09810570",
  1463 => x"b9d00807",
  1464 => x"9f2a7705",
  1465 => x"81175757",
  1466 => x"53537476",
  1467 => x"24893880",
  1468 => x"c0d40874",
  1469 => x"26d73872",
  1470 => x"b9d00c02",
  1471 => x"98050d04",
  1472 => x"02f0050d",
  1473 => x"b9cc0816",
  1474 => x"51adb62d",
  1475 => x"b9d00880",
  1476 => x"2e9c388b",
  1477 => x"53b9d008",
  1478 => x"52bec451",
  1479 => x"ad872d80",
  1480 => x"c1800854",
  1481 => x"73802e86",
  1482 => x"38bec451",
  1483 => x"732d0290",
  1484 => x"050d0402",
  1485 => x"dc050d80",
  1486 => x"705a5574",
  1487 => x"b9cc0825",
  1488 => x"b13880c0",
  1489 => x"d408752e",
  1490 => x"a9387851",
  1491 => x"a7a02db9",
  1492 => x"d0080981",
  1493 => x"0570b9d0",
  1494 => x"08079f2a",
  1495 => x"7605811b",
  1496 => x"5b565474",
  1497 => x"b9cc0825",
  1498 => x"893880c0",
  1499 => x"d4087926",
  1500 => x"d9388055",
  1501 => x"7880c0d4",
  1502 => x"082781d1",
  1503 => x"387851a7",
  1504 => x"a02db9d0",
  1505 => x"08802e81",
  1506 => x"a538b9d0",
  1507 => x"088b0580",
  1508 => x"f52d7084",
  1509 => x"2a708106",
  1510 => x"77107884",
  1511 => x"2bbec40b",
  1512 => x"80f52d5c",
  1513 => x"5c535155",
  1514 => x"5673802e",
  1515 => x"80c83874",
  1516 => x"16822bb0",
  1517 => x"f10bb8a0",
  1518 => x"120c5477",
  1519 => x"75311080",
  1520 => x"c1841155",
  1521 => x"56907470",
  1522 => x"81055681",
  1523 => x"b72da074",
  1524 => x"81b72d76",
  1525 => x"81ff0681",
  1526 => x"16585473",
  1527 => x"802e8938",
  1528 => x"9c53bec4",
  1529 => x"52afee04",
  1530 => x"8b53b9d0",
  1531 => x"085280c1",
  1532 => x"861651b0",
  1533 => x"a6047416",
  1534 => x"822bae80",
  1535 => x"0bb8a012",
  1536 => x"0c547681",
  1537 => x"ff068116",
  1538 => x"58547380",
  1539 => x"2e89389c",
  1540 => x"53bec452",
  1541 => x"b09d048b",
  1542 => x"53b9d008",
  1543 => x"52777531",
  1544 => x"1080c184",
  1545 => x"05517655",
  1546 => x"ad872db0",
  1547 => x"c2047490",
  1548 => x"29753170",
  1549 => x"1080c184",
  1550 => x"055154b9",
  1551 => x"d0087481",
  1552 => x"b72d8119",
  1553 => x"59748b24",
  1554 => x"a338aef4",
  1555 => x"04749029",
  1556 => x"75317010",
  1557 => x"80c18405",
  1558 => x"8c773157",
  1559 => x"51548074",
  1560 => x"81b72d9e",
  1561 => x"14ff1656",
  1562 => x"5474f338",
  1563 => x"02a4050d",
  1564 => x"0402fc05",
  1565 => x"0db9cc08",
  1566 => x"1351adb6",
  1567 => x"2db9d008",
  1568 => x"802e8838",
  1569 => x"b9d00851",
  1570 => x"9fcb2d80",
  1571 => x"0bb9cc0c",
  1572 => x"aeb32d8e",
  1573 => x"a82d0284",
  1574 => x"050d0402",
  1575 => x"fc050d72",
  1576 => x"5170fd2e",
  1577 => x"ad3870fd",
  1578 => x"248a3870",
  1579 => x"fc2e80c4",
  1580 => x"38b1fc04",
  1581 => x"70fe2eb1",
  1582 => x"3870ff2e",
  1583 => x"098106bc",
  1584 => x"38b9cc08",
  1585 => x"5170802e",
  1586 => x"b338ff11",
  1587 => x"b9cc0cb1",
  1588 => x"fc04b9cc",
  1589 => x"08f00570",
  1590 => x"b9cc0c51",
  1591 => x"7080259c",
  1592 => x"38800bb9",
  1593 => x"cc0cb1fc",
  1594 => x"04b9cc08",
  1595 => x"8105b9cc",
  1596 => x"0cb1fc04",
  1597 => x"b9cc0890",
  1598 => x"05b9cc0c",
  1599 => x"aeb32d8e",
  1600 => x"a82d0284",
  1601 => x"050d0402",
  1602 => x"fc050d80",
  1603 => x"0bb9cc0c",
  1604 => x"aeb32d8d",
  1605 => x"ad2db9d0",
  1606 => x"08b9bc0c",
  1607 => x"b898518f",
  1608 => x"c32d0284",
  1609 => x"050d0471",
  1610 => x"80c1800c",
  1611 => x"04000000",
  1612 => x"00ffffff",
  1613 => x"ff00ffff",
  1614 => x"ffff00ff",
  1615 => x"ffffff00",
  1616 => x"52657365",
  1617 => x"74000000",
  1618 => x"52474220",
  1619 => x"5363616c",
  1620 => x"696e6720",
  1621 => x"10000000",
  1622 => x"5363616e",
  1623 => x"6c696e65",
  1624 => x"73000000",
  1625 => x"416e696d",
  1626 => x"61746500",
  1627 => x"4c6f6164",
  1628 => x"20696d61",
  1629 => x"67652010",
  1630 => x"00000000",
  1631 => x"45786974",
  1632 => x"00000000",
  1633 => x"54657374",
  1634 => x"20706174",
  1635 => x"7465726e",
  1636 => x"20310000",
  1637 => x"54657374",
  1638 => x"20706174",
  1639 => x"7465726e",
  1640 => x"20320000",
  1641 => x"54657374",
  1642 => x"20706174",
  1643 => x"7465726e",
  1644 => x"20330000",
  1645 => x"54657374",
  1646 => x"20706174",
  1647 => x"7465726e",
  1648 => x"20340000",
  1649 => x"52656400",
  1650 => x"47726565",
  1651 => x"6e000000",
  1652 => x"426c7565",
  1653 => x"00000000",
  1654 => x"496e6974",
  1655 => x"69616c20",
  1656 => x"524f4d20",
  1657 => x"6c6f6164",
  1658 => x"696e6720",
  1659 => x"6661696c",
  1660 => x"65640000",
  1661 => x"4f4b0000",
  1662 => x"496e6974",
  1663 => x"69616c69",
  1664 => x"7a696e67",
  1665 => x"20534420",
  1666 => x"63617264",
  1667 => x"0a000000",
  1668 => x"4c6f6164",
  1669 => x"696e6720",
  1670 => x"696e6974",
  1671 => x"69616c20",
  1672 => x"524f4d2e",
  1673 => x"2e2e0a00",
  1674 => x"50494331",
  1675 => x"20202020",
  1676 => x"52415700",
  1677 => x"43617264",
  1678 => x"20696e69",
  1679 => x"74206661",
  1680 => x"696c6564",
  1681 => x"0a000000",
  1682 => x"16200000",
  1683 => x"14200000",
  1684 => x"15200000",
  1685 => x"53444843",
  1686 => x"20657272",
  1687 => x"6f72210a",
  1688 => x"00000000",
  1689 => x"53442069",
  1690 => x"6e69742e",
  1691 => x"2e2e0a00",
  1692 => x"53442063",
  1693 => x"61726420",
  1694 => x"72657365",
  1695 => x"74206661",
  1696 => x"696c6564",
  1697 => x"210a0000",
  1698 => x"57726974",
  1699 => x"65206661",
  1700 => x"696c6564",
  1701 => x"0a000000",
  1702 => x"52656164",
  1703 => x"20666169",
  1704 => x"6c65640a",
  1705 => x"00000000",
  1706 => x"4d425220",
  1707 => x"6661696c",
  1708 => x"0a000000",
  1709 => x"46415431",
  1710 => x"36202020",
  1711 => x"00000000",
  1712 => x"46415433",
  1713 => x"32202020",
  1714 => x"00000000",
  1715 => x"4e6f2070",
  1716 => x"61727469",
  1717 => x"74696f6e",
  1718 => x"20736967",
  1719 => x"0a000000",
  1720 => x"42616420",
  1721 => x"70617274",
  1722 => x"0a000000",
  1723 => x"4261636b",
  1724 => x"00000000",
  1725 => x"00000002",
  1726 => x"00000002",
  1727 => x"00001940",
  1728 => x"00000352",
  1729 => x"00000003",
  1730 => x"00001b58",
  1731 => x"00000004",
  1732 => x"00000004",
  1733 => x"00001948",
  1734 => x"00001b68",
  1735 => x"00000001",
  1736 => x"00001958",
  1737 => x"00000000",
  1738 => x"00000002",
  1739 => x"00001964",
  1740 => x"00000324",
  1741 => x"00000002",
  1742 => x"0000196c",
  1743 => x"00001907",
  1744 => x"00000002",
  1745 => x"0000197c",
  1746 => x"000006c7",
  1747 => x"00000000",
  1748 => x"00000000",
  1749 => x"00000000",
  1750 => x"00001984",
  1751 => x"00001994",
  1752 => x"000019a4",
  1753 => x"000019b4",
  1754 => x"00000005",
  1755 => x"000019c4",
  1756 => x"00000010",
  1757 => x"00000005",
  1758 => x"000019c8",
  1759 => x"00000010",
  1760 => x"00000005",
  1761 => x"000019d0",
  1762 => x"00000010",
  1763 => x"00000004",
  1764 => x"0000197c",
  1765 => x"00001af8",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000004",
  1770 => x"000019d8",
  1771 => x"00001ba4",
  1772 => x"00000004",
  1773 => x"000019f4",
  1774 => x"00001af8",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"00000000",
  1795 => x"00000000",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"00000002",
  1799 => x"00002084",
  1800 => x"00001700",
  1801 => x"00000002",
  1802 => x"000020a2",
  1803 => x"00001700",
  1804 => x"00000002",
  1805 => x"000020c0",
  1806 => x"00001700",
  1807 => x"00000002",
  1808 => x"000020de",
  1809 => x"00001700",
  1810 => x"00000002",
  1811 => x"000020fc",
  1812 => x"00001700",
  1813 => x"00000002",
  1814 => x"0000211a",
  1815 => x"00001700",
  1816 => x"00000002",
  1817 => x"00002138",
  1818 => x"00001700",
  1819 => x"00000002",
  1820 => x"00002156",
  1821 => x"00001700",
  1822 => x"00000002",
  1823 => x"00002174",
  1824 => x"00001700",
  1825 => x"00000002",
  1826 => x"00002192",
  1827 => x"00001700",
  1828 => x"00000002",
  1829 => x"000021b0",
  1830 => x"00001700",
  1831 => x"00000002",
  1832 => x"000021ce",
  1833 => x"00001700",
  1834 => x"00000002",
  1835 => x"000021ec",
  1836 => x"00001700",
  1837 => x"00000004",
  1838 => x"00001aec",
  1839 => x"00000000",
  1840 => x"00000000",
  1841 => x"00000000",
  1842 => x"0000189b",
  1843 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

