-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0b98",
     9 => x"c4080b0b",
    10 => x"0b98c808",
    11 => x"0b0b0b98",
    12 => x"cc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"98cc0c0b",
    16 => x"0b0b98c8",
    17 => x"0c0b0b0b",
    18 => x"98c40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0b95c4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"98c47099",
    57 => x"a8278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"85ec0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"98d40c9f",
    65 => x"0b98d80c",
    66 => x"a0717081",
    67 => x"05533498",
    68 => x"d808ff05",
    69 => x"98d80c98",
    70 => x"d8088025",
    71 => x"eb3898d4",
    72 => x"08ff0598",
    73 => x"d40c98d4",
    74 => x"088025d7",
    75 => x"38800b98",
    76 => x"d80c800b",
    77 => x"98d40c02",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"98d40825",
    97 => x"8f3882bc",
    98 => x"2d98d408",
    99 => x"ff0598d4",
   100 => x"0c82fe04",
   101 => x"98d40898",
   102 => x"d8085351",
   103 => x"728a2e09",
   104 => x"8106b738",
   105 => x"7151719f",
   106 => x"24a03898",
   107 => x"d408a029",
   108 => x"11f88011",
   109 => x"5151a071",
   110 => x"3498d808",
   111 => x"810598d8",
   112 => x"0c98d808",
   113 => x"519f7125",
   114 => x"e238800b",
   115 => x"98d80c98",
   116 => x"d4088105",
   117 => x"98d40c83",
   118 => x"ee0470a0",
   119 => x"2912f880",
   120 => x"11515172",
   121 => x"713498d8",
   122 => x"08810598",
   123 => x"d80c98d8",
   124 => x"08a02e09",
   125 => x"81068e38",
   126 => x"800b98d8",
   127 => x"0c98d408",
   128 => x"810598d4",
   129 => x"0c028c05",
   130 => x"0d0402ec",
   131 => x"050d800b",
   132 => x"98dc0cf6",
   133 => x"8c08f690",
   134 => x"0871882c",
   135 => x"565481ff",
   136 => x"06527372",
   137 => x"25883871",
   138 => x"54820b98",
   139 => x"dc0c7288",
   140 => x"2c7381ff",
   141 => x"06545574",
   142 => x"73258b38",
   143 => x"7298dc08",
   144 => x"840798dc",
   145 => x"0c557384",
   146 => x"2b86a071",
   147 => x"25837131",
   148 => x"700b0b0b",
   149 => x"96e00c81",
   150 => x"712bff05",
   151 => x"f6880cfe",
   152 => x"cc13ff12",
   153 => x"2c788829",
   154 => x"ff940570",
   155 => x"812c98dc",
   156 => x"08525852",
   157 => x"55515254",
   158 => x"76802e85",
   159 => x"38708107",
   160 => x"5170f694",
   161 => x"0c710981",
   162 => x"05f6800c",
   163 => x"72098105",
   164 => x"f6840c02",
   165 => x"94050d04",
   166 => x"02f4050d",
   167 => x"74537270",
   168 => x"81055480",
   169 => x"f52d5271",
   170 => x"802e8938",
   171 => x"715182f8",
   172 => x"2d859e04",
   173 => x"810b98c4",
   174 => x"0c028c05",
   175 => x"0d0402fc",
   176 => x"050d8acd",
   177 => x"2d80518a",
   178 => x"872d8a87",
   179 => x"2d8a872d",
   180 => x"8a872d70",
   181 => x"f00c70f4",
   182 => x"0c70f80c",
   183 => x"81115190",
   184 => x"7125e438",
   185 => x"8aba2d02",
   186 => x"84050d04",
   187 => x"02f4050d",
   188 => x"8aa22d86",
   189 => x"f12d81f7",
   190 => x"2d97a051",
   191 => x"8cab2d83",
   192 => x"528a872d",
   193 => x"8151848a",
   194 => x"2dff1252",
   195 => x"718025f1",
   196 => x"38880b96",
   197 => x"ec0b81b7",
   198 => x"2d880b96",
   199 => x"f80b81b7",
   200 => x"2d880b97",
   201 => x"840b81b7",
   202 => x"2d8aba2d",
   203 => x"86fd2d8c",
   204 => x"bb2d97a8",
   205 => x"0b80f52d",
   206 => x"998c0881",
   207 => x"06535371",
   208 => x"802e8538",
   209 => x"72840753",
   210 => x"72fc0c96",
   211 => x"ec0b80f5",
   212 => x"2df00c96",
   213 => x"f80b80f5",
   214 => x"2df40c97",
   215 => x"840b80f5",
   216 => x"2df80c86",
   217 => x"ac047198",
   218 => x"0c04ffb0",
   219 => x"0898c40c",
   220 => x"04810bff",
   221 => x"b00c0480",
   222 => x"0bffb00c",
   223 => x"0402f405",
   224 => x"0d87ff04",
   225 => x"98c40881",
   226 => x"f02e0981",
   227 => x"06893881",
   228 => x"0b98b80c",
   229 => x"87ff0498",
   230 => x"c40881e0",
   231 => x"2e098106",
   232 => x"8938810b",
   233 => x"98bc0c87",
   234 => x"ff0498c4",
   235 => x"085298bc",
   236 => x"08802e88",
   237 => x"3898c408",
   238 => x"81800552",
   239 => x"71842c72",
   240 => x"8f065353",
   241 => x"98b80880",
   242 => x"2e993872",
   243 => x"842997f8",
   244 => x"05721381",
   245 => x"712b7009",
   246 => x"73080673",
   247 => x"0c515353",
   248 => x"87f50472",
   249 => x"842997f8",
   250 => x"05721383",
   251 => x"712b7208",
   252 => x"07720c53",
   253 => x"53800b98",
   254 => x"bc0c800b",
   255 => x"98b80c98",
   256 => x"e0518980",
   257 => x"2d98c408",
   258 => x"ff24fef8",
   259 => x"38800b98",
   260 => x"c40c028c",
   261 => x"050d0402",
   262 => x"f8050d97",
   263 => x"f8528f51",
   264 => x"80727084",
   265 => x"05540cff",
   266 => x"11517080",
   267 => x"25f23802",
   268 => x"88050d04",
   269 => x"02f0050d",
   270 => x"755186f7",
   271 => x"2d70822c",
   272 => x"fc0697f8",
   273 => x"1172109e",
   274 => x"06710870",
   275 => x"722a7083",
   276 => x"0682742b",
   277 => x"70097406",
   278 => x"760c5451",
   279 => x"56575351",
   280 => x"5386f12d",
   281 => x"7198c40c",
   282 => x"0290050d",
   283 => x"0402fc05",
   284 => x"0d725180",
   285 => x"710c800b",
   286 => x"84120c02",
   287 => x"84050d04",
   288 => x"02f0050d",
   289 => x"75700884",
   290 => x"12085353",
   291 => x"53ff5471",
   292 => x"712ea838",
   293 => x"86f72d84",
   294 => x"13087084",
   295 => x"29148811",
   296 => x"70087081",
   297 => x"ff068418",
   298 => x"08811187",
   299 => x"06841a0c",
   300 => x"53515551",
   301 => x"515186f1",
   302 => x"2d715473",
   303 => x"98c40c02",
   304 => x"90050d04",
   305 => x"02f8050d",
   306 => x"86f72de0",
   307 => x"08708b2a",
   308 => x"70810651",
   309 => x"52527080",
   310 => x"2e9d3898",
   311 => x"e0087084",
   312 => x"2998e805",
   313 => x"7381ff06",
   314 => x"710c5151",
   315 => x"98e00881",
   316 => x"11870698",
   317 => x"e00c5180",
   318 => x"0b99880c",
   319 => x"86ea2d86",
   320 => x"f12d0288",
   321 => x"050d0402",
   322 => x"fc050d86",
   323 => x"f72d810b",
   324 => x"99880c86",
   325 => x"f12d9988",
   326 => x"085170fa",
   327 => x"38028405",
   328 => x"0d0402fc",
   329 => x"050d98e0",
   330 => x"5188ed2d",
   331 => x"88972d89",
   332 => x"c45186e6",
   333 => x"2d028405",
   334 => x"0d0402fc",
   335 => x"050d810b",
   336 => x"98c00c81",
   337 => x"51848a2d",
   338 => x"0284050d",
   339 => x"0402fc05",
   340 => x"0d800b98",
   341 => x"c00c8051",
   342 => x"848a2d02",
   343 => x"84050d04",
   344 => x"02ec050d",
   345 => x"76548052",
   346 => x"870b8815",
   347 => x"80f52d56",
   348 => x"53747224",
   349 => x"8338a053",
   350 => x"725182f8",
   351 => x"2d81128b",
   352 => x"1580f52d",
   353 => x"54527272",
   354 => x"25de3802",
   355 => x"94050d04",
   356 => x"02f0050d",
   357 => x"99980854",
   358 => x"81f72d80",
   359 => x"0b999c0c",
   360 => x"7308802e",
   361 => x"81803882",
   362 => x"0b98d80c",
   363 => x"999c088f",
   364 => x"0698d40c",
   365 => x"73085271",
   366 => x"832e9638",
   367 => x"71832689",
   368 => x"3871812e",
   369 => x"af388c91",
   370 => x"0471852e",
   371 => x"9f388c91",
   372 => x"04881480",
   373 => x"f52d8415",
   374 => x"0896d453",
   375 => x"54528598",
   376 => x"2d718429",
   377 => x"13700852",
   378 => x"528c9504",
   379 => x"73518ae0",
   380 => x"2d8c9104",
   381 => x"998c0888",
   382 => x"15082c70",
   383 => x"81065152",
   384 => x"71802e87",
   385 => x"3896d851",
   386 => x"8c8e0496",
   387 => x"dc518598",
   388 => x"2d841408",
   389 => x"5185982d",
   390 => x"999c0881",
   391 => x"05999c0c",
   392 => x"8c14548b",
   393 => x"a0040290",
   394 => x"050d0471",
   395 => x"99980c8b",
   396 => x"902d999c",
   397 => x"08ff0599",
   398 => x"a00c0402",
   399 => x"e8050d99",
   400 => x"980899a4",
   401 => x"08575580",
   402 => x"f85188b4",
   403 => x"2d98c408",
   404 => x"812a7081",
   405 => x"06515271",
   406 => x"9b388751",
   407 => x"88b42d98",
   408 => x"c408812a",
   409 => x"70810651",
   410 => x"5271802e",
   411 => x"b1388cf4",
   412 => x"0486fd2d",
   413 => x"875188b4",
   414 => x"2d98c408",
   415 => x"f4388d84",
   416 => x"0486fd2d",
   417 => x"80f85188",
   418 => x"b42d98c4",
   419 => x"08f33898",
   420 => x"c0088132",
   421 => x"7098c00c",
   422 => x"70525284",
   423 => x"8a2d800b",
   424 => x"99900c80",
   425 => x"0b99940c",
   426 => x"98c00882",
   427 => x"dd3880da",
   428 => x"5188b42d",
   429 => x"98c40880",
   430 => x"2e8a3899",
   431 => x"90088180",
   432 => x"0799900c",
   433 => x"80d95188",
   434 => x"b42d98c4",
   435 => x"08802e8a",
   436 => x"38999008",
   437 => x"80c00799",
   438 => x"900c8194",
   439 => x"5188b42d",
   440 => x"98c40880",
   441 => x"2e893899",
   442 => x"90089007",
   443 => x"99900c81",
   444 => x"915188b4",
   445 => x"2d98c408",
   446 => x"802e8938",
   447 => x"999008a0",
   448 => x"0799900c",
   449 => x"81f55188",
   450 => x"b42d98c4",
   451 => x"08802e89",
   452 => x"38999008",
   453 => x"81079990",
   454 => x"0c81f251",
   455 => x"88b42d98",
   456 => x"c408802e",
   457 => x"89389990",
   458 => x"08820799",
   459 => x"900c81eb",
   460 => x"5188b42d",
   461 => x"98c40880",
   462 => x"2e893899",
   463 => x"90088407",
   464 => x"99900c81",
   465 => x"f45188b4",
   466 => x"2d98c408",
   467 => x"802e8938",
   468 => x"99900888",
   469 => x"0799900c",
   470 => x"80d85188",
   471 => x"b42d98c4",
   472 => x"08802e8a",
   473 => x"38999408",
   474 => x"81800799",
   475 => x"940c9251",
   476 => x"88b42d98",
   477 => x"c408802e",
   478 => x"8a389994",
   479 => x"0880c007",
   480 => x"99940c94",
   481 => x"5188b42d",
   482 => x"98c40880",
   483 => x"2e893899",
   484 => x"94089007",
   485 => x"99940c91",
   486 => x"5188b42d",
   487 => x"98c40880",
   488 => x"2e893899",
   489 => x"9408a007",
   490 => x"99940c9d",
   491 => x"5188b42d",
   492 => x"98c40880",
   493 => x"2e893899",
   494 => x"94088107",
   495 => x"99940c9b",
   496 => x"5188b42d",
   497 => x"98c40880",
   498 => x"2e893899",
   499 => x"94088207",
   500 => x"99940c9c",
   501 => x"5188b42d",
   502 => x"98c40880",
   503 => x"2e893899",
   504 => x"94088407",
   505 => x"99940ca3",
   506 => x"5188b42d",
   507 => x"98c40880",
   508 => x"2e893899",
   509 => x"94088807",
   510 => x"99940c81",
   511 => x"fd5188b4",
   512 => x"2d81fa51",
   513 => x"88b42d95",
   514 => x"bb0481f5",
   515 => x"5188b42d",
   516 => x"98c40881",
   517 => x"2a708106",
   518 => x"51527180",
   519 => x"2eaf3899",
   520 => x"a0085271",
   521 => x"802e8938",
   522 => x"ff1299a0",
   523 => x"0c90cd04",
   524 => x"999c0810",
   525 => x"999c0805",
   526 => x"70842916",
   527 => x"51528812",
   528 => x"08802e89",
   529 => x"38ff5188",
   530 => x"12085271",
   531 => x"2d81f251",
   532 => x"88b42d98",
   533 => x"c408812a",
   534 => x"70810651",
   535 => x"5271802e",
   536 => x"b138999c",
   537 => x"08ff1199",
   538 => x"a0085653",
   539 => x"53737225",
   540 => x"89388114",
   541 => x"99a00c91",
   542 => x"92047210",
   543 => x"13708429",
   544 => x"16515288",
   545 => x"1208802e",
   546 => x"8938fe51",
   547 => x"88120852",
   548 => x"712d81fd",
   549 => x"5188b42d",
   550 => x"98c40881",
   551 => x"2a708106",
   552 => x"51527180",
   553 => x"2ead3899",
   554 => x"a008802e",
   555 => x"8938800b",
   556 => x"99a00c91",
   557 => x"d304999c",
   558 => x"0810999c",
   559 => x"08057084",
   560 => x"29165152",
   561 => x"88120880",
   562 => x"2e8938fd",
   563 => x"51881208",
   564 => x"52712d81",
   565 => x"fa5188b4",
   566 => x"2d98c408",
   567 => x"812a7081",
   568 => x"06515271",
   569 => x"802eae38",
   570 => x"999c08ff",
   571 => x"11545299",
   572 => x"a0087325",
   573 => x"88387299",
   574 => x"a00c9295",
   575 => x"04711012",
   576 => x"70842916",
   577 => x"51528812",
   578 => x"08802e89",
   579 => x"38fc5188",
   580 => x"12085271",
   581 => x"2d99a008",
   582 => x"70535473",
   583 => x"802e8a38",
   584 => x"8c15ff15",
   585 => x"5555929b",
   586 => x"04820b98",
   587 => x"d80c718f",
   588 => x"0698d40c",
   589 => x"81eb5188",
   590 => x"b42d98c4",
   591 => x"08812a70",
   592 => x"81065152",
   593 => x"71802ead",
   594 => x"38740885",
   595 => x"2e098106",
   596 => x"a4388815",
   597 => x"80f52dff",
   598 => x"05527188",
   599 => x"1681b72d",
   600 => x"71982b52",
   601 => x"71802588",
   602 => x"38800b88",
   603 => x"1681b72d",
   604 => x"74518ae0",
   605 => x"2d81f451",
   606 => x"88b42d98",
   607 => x"c408812a",
   608 => x"70810651",
   609 => x"5271802e",
   610 => x"b3387408",
   611 => x"852e0981",
   612 => x"06aa3888",
   613 => x"1580f52d",
   614 => x"81055271",
   615 => x"881681b7",
   616 => x"2d7181ff",
   617 => x"068b1680",
   618 => x"f52d5452",
   619 => x"72722787",
   620 => x"38728816",
   621 => x"81b72d74",
   622 => x"518ae02d",
   623 => x"80da5188",
   624 => x"b42d98c4",
   625 => x"08812a70",
   626 => x"81065152",
   627 => x"71802e81",
   628 => x"a6389998",
   629 => x"0899a008",
   630 => x"55537380",
   631 => x"2e8a388c",
   632 => x"13ff1555",
   633 => x"5393da04",
   634 => x"72085271",
   635 => x"822ea638",
   636 => x"71822689",
   637 => x"3871812e",
   638 => x"a93894f7",
   639 => x"0471832e",
   640 => x"b1387184",
   641 => x"2e098106",
   642 => x"80ed3888",
   643 => x"1308518c",
   644 => x"ab2d94f7",
   645 => x"0499a008",
   646 => x"51881308",
   647 => x"52712d94",
   648 => x"f704810b",
   649 => x"8814082b",
   650 => x"998c0832",
   651 => x"998c0c94",
   652 => x"cd048813",
   653 => x"80f52d81",
   654 => x"058b1480",
   655 => x"f52d5354",
   656 => x"71742483",
   657 => x"38805473",
   658 => x"881481b7",
   659 => x"2d8b902d",
   660 => x"94f70475",
   661 => x"08802ea2",
   662 => x"38750851",
   663 => x"88b42d98",
   664 => x"c4088106",
   665 => x"5271802e",
   666 => x"8b3899a0",
   667 => x"08518416",
   668 => x"0852712d",
   669 => x"88165675",
   670 => x"da388054",
   671 => x"800b98d8",
   672 => x"0c738f06",
   673 => x"98d40ca0",
   674 => x"527399a0",
   675 => x"082e0981",
   676 => x"06983899",
   677 => x"9c08ff05",
   678 => x"74327009",
   679 => x"81057072",
   680 => x"079f2a91",
   681 => x"71315151",
   682 => x"53537151",
   683 => x"82f82d81",
   684 => x"14548e74",
   685 => x"25c63898",
   686 => x"c0085271",
   687 => x"98c40c02",
   688 => x"98050d04",
   689 => x"00ffffff",
   690 => x"ff00ffff",
   691 => x"ffff00ff",
   692 => x"ffffff00",
   693 => x"52656400",
   694 => x"47726565",
   695 => x"6e000000",
   696 => x"426c7565",
   697 => x"00000000",
   698 => x"45786974",
   699 => x"00000000",
   700 => x"52474220",
   701 => x"5363616c",
   702 => x"696e6720",
   703 => x"10000000",
   704 => x"5363616e",
   705 => x"6c696e65",
   706 => x"73000000",
   707 => x"416e696d",
   708 => x"61746500",
   709 => x"54657374",
   710 => x"20706174",
   711 => x"7465726e",
   712 => x"20310000",
   713 => x"54657374",
   714 => x"20706174",
   715 => x"7465726e",
   716 => x"20320000",
   717 => x"54657374",
   718 => x"20706174",
   719 => x"7465726e",
   720 => x"20330000",
   721 => x"54657374",
   722 => x"20706174",
   723 => x"7465726e",
   724 => x"20340000",
   725 => x"16200000",
   726 => x"14200000",
   727 => x"15200000",
   728 => x"00000002",
   729 => x"00000005",
   730 => x"00000ad4",
   731 => x"00000010",
   732 => x"00000005",
   733 => x"00000ad8",
   734 => x"00000010",
   735 => x"00000005",
   736 => x"00000ae0",
   737 => x"00000010",
   738 => x"00000004",
   739 => x"00000ae8",
   740 => x"00000ba0",
   741 => x"00000000",
   742 => x"00000000",
   743 => x"00000000",
   744 => x"00000003",
   745 => x"00000be8",
   746 => x"00000004",
   747 => x"00000004",
   748 => x"00000af0",
   749 => x"00000b64",
   750 => x"00000001",
   751 => x"00000b00",
   752 => x"00000000",
   753 => x"00000002",
   754 => x"00000b0c",
   755 => x"000002be",
   756 => x"00000002",
   757 => x"00000ae8",
   758 => x"0000054d",
   759 => x"00000000",
   760 => x"00000000",
   761 => x"00000000",
   762 => x"00000b14",
   763 => x"00000b24",
   764 => x"00000b34",
   765 => x"00000b44",
   766 => x"00000000",
   767 => x"00000000",
   768 => x"00000000",
   769 => x"00000000",
   770 => x"00000000",
   771 => x"00000000",
   772 => x"00000000",
   773 => x"00000000",
   774 => x"00000000",
   775 => x"00000000",
   776 => x"00000000",
   777 => x"00000000",
   778 => x"00000000",
   779 => x"00000000",
   780 => x"00000000",
   781 => x"00000000",
   782 => x"00000000",
   783 => x"00000000",
   784 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

