-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb9",
     9 => x"8c080b0b",
    10 => x"0bb99008",
    11 => x"0b0b0bb9",
    12 => x"94080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b9940c0b",
    16 => x"0b0bb990",
    17 => x"0c0b0b0b",
    18 => x"b98c0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb1f8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b98c7080",
    57 => x"c3c8278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"51888804",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb99c0c",
    65 => x"9f0bb9a0",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b9a008ff",
    69 => x"05b9a00c",
    70 => x"b9a00880",
    71 => x"25eb38b9",
    72 => x"9c08ff05",
    73 => x"b99c0cb9",
    74 => x"9c088025",
    75 => x"d738800b",
    76 => x"b9a00c80",
    77 => x"0bb99c0c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb99c08",
    97 => x"258f3882",
    98 => x"bd2db99c",
    99 => x"08ff05b9",
   100 => x"9c0c82ff",
   101 => x"04b99c08",
   102 => x"b9a00853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b99c08a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b9a0",
   111 => x"088105b9",
   112 => x"a00cb9a0",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb9a00c",
   116 => x"b99c0881",
   117 => x"05b99c0c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b9",
   122 => x"a0088105",
   123 => x"b9a00cb9",
   124 => x"a008a02e",
   125 => x"0981068e",
   126 => x"38800bb9",
   127 => x"a00cb99c",
   128 => x"088105b9",
   129 => x"9c0c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb9a4",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb9a40c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b9",
   169 => x"a4088407",
   170 => x"b9a40c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb5b0",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfecc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b9a40852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b98c0c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"8dab2d80",
   203 => x"518cde2d",
   204 => x"8cde2d8c",
   205 => x"de2d8cde",
   206 => x"2d70f00c",
   207 => x"70f40c70",
   208 => x"f80c8111",
   209 => x"51907125",
   210 => x"e4388d98",
   211 => x"2d028405",
   212 => x"0d0402fc",
   213 => x"050dec51",
   214 => x"83710c82",
   215 => x"710c0284",
   216 => x"050d0402",
   217 => x"dc050d80",
   218 => x"59810bec",
   219 => x"0c840bec",
   220 => x"0c7a52b9",
   221 => x"a851a99d",
   222 => x"2db98c08",
   223 => x"792e80f9",
   224 => x"38b9ac08",
   225 => x"79ff1256",
   226 => x"59567379",
   227 => x"2e8b3881",
   228 => x"1874812a",
   229 => x"555873f7",
   230 => x"38f71858",
   231 => x"81598076",
   232 => x"2580d038",
   233 => x"77527351",
   234 => x"848b2dba",
   235 => x"8052b9a8",
   236 => x"51abdc2d",
   237 => x"b98c0880",
   238 => x"2e9a38ba",
   239 => x"805783fc",
   240 => x"55767084",
   241 => x"055808e8",
   242 => x"0cfc1555",
   243 => x"748025f1",
   244 => x"3887db04",
   245 => x"b98c0859",
   246 => x"848056b9",
   247 => x"a851abae",
   248 => x"2dfc8016",
   249 => x"81155556",
   250 => x"758024ff",
   251 => x"b7387880",
   252 => x"2e8738b5",
   253 => x"b45187fc",
   254 => x"04b6e051",
   255 => x"8fa72d78",
   256 => x"b98c0c02",
   257 => x"a4050d04",
   258 => x"02f4050d",
   259 => x"810bec0c",
   260 => x"8cf92d89",
   261 => x"c82d81f8",
   262 => x"2d83528c",
   263 => x"de2d8151",
   264 => x"84f02dff",
   265 => x"12527180",
   266 => x"25f13888",
   267 => x"0bb6ac0b",
   268 => x"81b72d88",
   269 => x"0bb6b80b",
   270 => x"81b72d88",
   271 => x"0bb6c40b",
   272 => x"81b72d84",
   273 => x"0bec0cb3",
   274 => x"c05185fe",
   275 => x"2da09c2d",
   276 => x"b98c0880",
   277 => x"2e80dc38",
   278 => x"b3d85185",
   279 => x"fe2db3f0",
   280 => x"5186e32d",
   281 => x"86e351b1",
   282 => x"f12d8d98",
   283 => x"2d89d42d",
   284 => x"8fb72db5",
   285 => x"c80b80f5",
   286 => x"2db9e008",
   287 => x"81065353",
   288 => x"71802e85",
   289 => x"38728407",
   290 => x"5372fc0c",
   291 => x"b6ac0b80",
   292 => x"f52df00c",
   293 => x"b6b80b80",
   294 => x"f52df40c",
   295 => x"b6c40b80",
   296 => x"f52df80c",
   297 => x"8652b98c",
   298 => x"08833884",
   299 => x"5271ec0c",
   300 => x"88ed0480",
   301 => x"0bb98c0c",
   302 => x"028c050d",
   303 => x"0471980c",
   304 => x"04ffb008",
   305 => x"b98c0c04",
   306 => x"810bffb0",
   307 => x"0c04800b",
   308 => x"ffb00c04",
   309 => x"02f4050d",
   310 => x"8ad604b9",
   311 => x"8c0881f0",
   312 => x"2e098106",
   313 => x"8938810b",
   314 => x"b7c40c8a",
   315 => x"d604b98c",
   316 => x"0881e02e",
   317 => x"09810689",
   318 => x"38810bb7",
   319 => x"c80c8ad6",
   320 => x"04b98c08",
   321 => x"52b7c808",
   322 => x"802e8838",
   323 => x"b98c0881",
   324 => x"80055271",
   325 => x"842c728f",
   326 => x"065353b7",
   327 => x"c408802e",
   328 => x"99387284",
   329 => x"29b78405",
   330 => x"72138171",
   331 => x"2b700973",
   332 => x"0806730c",
   333 => x"5153538a",
   334 => x"cc047284",
   335 => x"29b78405",
   336 => x"72138371",
   337 => x"2b720807",
   338 => x"720c5353",
   339 => x"800bb7c8",
   340 => x"0c800bb7",
   341 => x"c40cb9b4",
   342 => x"518bd72d",
   343 => x"b98c08ff",
   344 => x"24fef838",
   345 => x"800bb98c",
   346 => x"0c028c05",
   347 => x"0d0402f8",
   348 => x"050db784",
   349 => x"528f5180",
   350 => x"72708405",
   351 => x"540cff11",
   352 => x"51708025",
   353 => x"f2380288",
   354 => x"050d0402",
   355 => x"f0050d75",
   356 => x"5189ce2d",
   357 => x"70822cfc",
   358 => x"06b78411",
   359 => x"72109e06",
   360 => x"71087072",
   361 => x"2a708306",
   362 => x"82742b70",
   363 => x"09740676",
   364 => x"0c545156",
   365 => x"57535153",
   366 => x"89c82d71",
   367 => x"b98c0c02",
   368 => x"90050d04",
   369 => x"02fc050d",
   370 => x"72518071",
   371 => x"0c800b84",
   372 => x"120c0284",
   373 => x"050d0402",
   374 => x"f0050d75",
   375 => x"70088412",
   376 => x"08535353",
   377 => x"ff547171",
   378 => x"2ea83889",
   379 => x"ce2d8413",
   380 => x"08708429",
   381 => x"14881170",
   382 => x"087081ff",
   383 => x"06841808",
   384 => x"81118706",
   385 => x"841a0c53",
   386 => x"51555151",
   387 => x"5189c82d",
   388 => x"715473b9",
   389 => x"8c0c0290",
   390 => x"050d0402",
   391 => x"f8050d89",
   392 => x"ce2de008",
   393 => x"708b2a70",
   394 => x"81065152",
   395 => x"5270802e",
   396 => x"9d38b9b4",
   397 => x"08708429",
   398 => x"b9bc0573",
   399 => x"81ff0671",
   400 => x"0c5151b9",
   401 => x"b4088111",
   402 => x"8706b9b4",
   403 => x"0c51800b",
   404 => x"b9dc0c89",
   405 => x"c12d89c8",
   406 => x"2d028805",
   407 => x"0d0402fc",
   408 => x"050d89ce",
   409 => x"2d810bb9",
   410 => x"dc0c89c8",
   411 => x"2db9dc08",
   412 => x"5170fa38",
   413 => x"0284050d",
   414 => x"0402fc05",
   415 => x"0db9b451",
   416 => x"8bc42d8a",
   417 => x"ee2d8c9b",
   418 => x"5189bd2d",
   419 => x"0284050d",
   420 => x"04b9ec08",
   421 => x"b98c0c04",
   422 => x"02fc050d",
   423 => x"810bb7cc",
   424 => x"0c815184",
   425 => x"f02d0284",
   426 => x"050d0402",
   427 => x"fc050d8d",
   428 => x"b50489d4",
   429 => x"2d87518b",
   430 => x"8b2db98c",
   431 => x"08f43880",
   432 => x"da518b8b",
   433 => x"2db98c08",
   434 => x"e938b98c",
   435 => x"08b7cc0c",
   436 => x"b98c0851",
   437 => x"84f02d02",
   438 => x"84050d04",
   439 => x"02ec050d",
   440 => x"76548052",
   441 => x"870b8815",
   442 => x"80f52d56",
   443 => x"53747224",
   444 => x"8338a053",
   445 => x"725182f9",
   446 => x"2d81128b",
   447 => x"1580f52d",
   448 => x"54527272",
   449 => x"25de3802",
   450 => x"94050d04",
   451 => x"02f0050d",
   452 => x"b9ec0854",
   453 => x"81f82d80",
   454 => x"0bb9f00c",
   455 => x"7308802e",
   456 => x"81803882",
   457 => x"0bb9a00c",
   458 => x"b9f0088f",
   459 => x"06b99c0c",
   460 => x"73085271",
   461 => x"832e9638",
   462 => x"71832689",
   463 => x"3871812e",
   464 => x"af388f8d",
   465 => x"0471852e",
   466 => x"9f388f8d",
   467 => x"04881480",
   468 => x"f52d8415",
   469 => x"08b3fc53",
   470 => x"545285fe",
   471 => x"2d718429",
   472 => x"13700852",
   473 => x"528f9104",
   474 => x"73518ddc",
   475 => x"2d8f8d04",
   476 => x"b9e00888",
   477 => x"15082c70",
   478 => x"81065152",
   479 => x"71802e87",
   480 => x"38b48051",
   481 => x"8f8a04b4",
   482 => x"845185fe",
   483 => x"2d841408",
   484 => x"5185fe2d",
   485 => x"b9f00881",
   486 => x"05b9f00c",
   487 => x"8c14548e",
   488 => x"9c040290",
   489 => x"050d0471",
   490 => x"b9ec0c8e",
   491 => x"8c2db9f0",
   492 => x"08ff05b9",
   493 => x"f40c0402",
   494 => x"e8050db9",
   495 => x"ec08b9f8",
   496 => x"08575587",
   497 => x"518b8b2d",
   498 => x"b98c0881",
   499 => x"2a708106",
   500 => x"51527180",
   501 => x"2ea0388f",
   502 => x"dd0489d4",
   503 => x"2d87518b",
   504 => x"8b2db98c",
   505 => x"08f438b7",
   506 => x"cc088132",
   507 => x"70b7cc0c",
   508 => x"70525284",
   509 => x"f02d800b",
   510 => x"b9e40c80",
   511 => x"0bb9e80c",
   512 => x"b7cc0882",
   513 => x"dd3880da",
   514 => x"518b8b2d",
   515 => x"b98c0880",
   516 => x"2e8a38b9",
   517 => x"e4088180",
   518 => x"07b9e40c",
   519 => x"80d9518b",
   520 => x"8b2db98c",
   521 => x"08802e8a",
   522 => x"38b9e408",
   523 => x"80c007b9",
   524 => x"e40c8194",
   525 => x"518b8b2d",
   526 => x"b98c0880",
   527 => x"2e8938b9",
   528 => x"e4089007",
   529 => x"b9e40c81",
   530 => x"91518b8b",
   531 => x"2db98c08",
   532 => x"802e8938",
   533 => x"b9e408a0",
   534 => x"07b9e40c",
   535 => x"81f5518b",
   536 => x"8b2db98c",
   537 => x"08802e89",
   538 => x"38b9e408",
   539 => x"8107b9e4",
   540 => x"0c81f251",
   541 => x"8b8b2db9",
   542 => x"8c08802e",
   543 => x"8938b9e4",
   544 => x"088207b9",
   545 => x"e40c81eb",
   546 => x"518b8b2d",
   547 => x"b98c0880",
   548 => x"2e8938b9",
   549 => x"e4088407",
   550 => x"b9e40c81",
   551 => x"f4518b8b",
   552 => x"2db98c08",
   553 => x"802e8938",
   554 => x"b9e40888",
   555 => x"07b9e40c",
   556 => x"80d8518b",
   557 => x"8b2db98c",
   558 => x"08802e8a",
   559 => x"38b9e808",
   560 => x"818007b9",
   561 => x"e80c9251",
   562 => x"8b8b2db9",
   563 => x"8c08802e",
   564 => x"8a38b9e8",
   565 => x"0880c007",
   566 => x"b9e80c94",
   567 => x"518b8b2d",
   568 => x"b98c0880",
   569 => x"2e8938b9",
   570 => x"e8089007",
   571 => x"b9e80c91",
   572 => x"518b8b2d",
   573 => x"b98c0880",
   574 => x"2e8938b9",
   575 => x"e808a007",
   576 => x"b9e80c9d",
   577 => x"518b8b2d",
   578 => x"b98c0880",
   579 => x"2e8938b9",
   580 => x"e8088107",
   581 => x"b9e80c9b",
   582 => x"518b8b2d",
   583 => x"b98c0880",
   584 => x"2e8938b9",
   585 => x"e8088207",
   586 => x"b9e80c9c",
   587 => x"518b8b2d",
   588 => x"b98c0880",
   589 => x"2e8938b9",
   590 => x"e8088407",
   591 => x"b9e80ca3",
   592 => x"518b8b2d",
   593 => x"b98c0880",
   594 => x"2e8938b9",
   595 => x"e8088807",
   596 => x"b9e80c81",
   597 => x"fd518b8b",
   598 => x"2d81fa51",
   599 => x"8b8b2d98",
   600 => x"930481f5",
   601 => x"518b8b2d",
   602 => x"b98c0881",
   603 => x"2a708106",
   604 => x"51527180",
   605 => x"2eaf38b9",
   606 => x"f4085271",
   607 => x"802e8938",
   608 => x"ff12b9f4",
   609 => x"0c93a504",
   610 => x"b9f00810",
   611 => x"b9f00805",
   612 => x"70842916",
   613 => x"51528812",
   614 => x"08802e89",
   615 => x"38ff5188",
   616 => x"12085271",
   617 => x"2d81f251",
   618 => x"8b8b2db9",
   619 => x"8c08812a",
   620 => x"70810651",
   621 => x"5271802e",
   622 => x"b138b9f0",
   623 => x"08ff11b9",
   624 => x"f4085653",
   625 => x"53737225",
   626 => x"89388114",
   627 => x"b9f40c93",
   628 => x"ea047210",
   629 => x"13708429",
   630 => x"16515288",
   631 => x"1208802e",
   632 => x"8938fe51",
   633 => x"88120852",
   634 => x"712d81fd",
   635 => x"518b8b2d",
   636 => x"b98c0881",
   637 => x"2a708106",
   638 => x"51527180",
   639 => x"2ead38b9",
   640 => x"f408802e",
   641 => x"8938800b",
   642 => x"b9f40c94",
   643 => x"ab04b9f0",
   644 => x"0810b9f0",
   645 => x"08057084",
   646 => x"29165152",
   647 => x"88120880",
   648 => x"2e8938fd",
   649 => x"51881208",
   650 => x"52712d81",
   651 => x"fa518b8b",
   652 => x"2db98c08",
   653 => x"812a7081",
   654 => x"06515271",
   655 => x"802eae38",
   656 => x"b9f008ff",
   657 => x"115452b9",
   658 => x"f4087325",
   659 => x"883872b9",
   660 => x"f40c94ed",
   661 => x"04711012",
   662 => x"70842916",
   663 => x"51528812",
   664 => x"08802e89",
   665 => x"38fc5188",
   666 => x"12085271",
   667 => x"2db9f408",
   668 => x"70535473",
   669 => x"802e8a38",
   670 => x"8c15ff15",
   671 => x"555594f3",
   672 => x"04820bb9",
   673 => x"a00c718f",
   674 => x"06b99c0c",
   675 => x"81eb518b",
   676 => x"8b2db98c",
   677 => x"08812a70",
   678 => x"81065152",
   679 => x"71802ead",
   680 => x"38740885",
   681 => x"2e098106",
   682 => x"a4388815",
   683 => x"80f52dff",
   684 => x"05527188",
   685 => x"1681b72d",
   686 => x"71982b52",
   687 => x"71802588",
   688 => x"38800b88",
   689 => x"1681b72d",
   690 => x"74518ddc",
   691 => x"2d81f451",
   692 => x"8b8b2db9",
   693 => x"8c08812a",
   694 => x"70810651",
   695 => x"5271802e",
   696 => x"b3387408",
   697 => x"852e0981",
   698 => x"06aa3888",
   699 => x"1580f52d",
   700 => x"81055271",
   701 => x"881681b7",
   702 => x"2d7181ff",
   703 => x"068b1680",
   704 => x"f52d5452",
   705 => x"72722787",
   706 => x"38728816",
   707 => x"81b72d74",
   708 => x"518ddc2d",
   709 => x"80da518b",
   710 => x"8b2db98c",
   711 => x"08812a70",
   712 => x"81065152",
   713 => x"71802e81",
   714 => x"a638b9ec",
   715 => x"08b9f408",
   716 => x"55537380",
   717 => x"2e8a388c",
   718 => x"13ff1555",
   719 => x"5396b204",
   720 => x"72085271",
   721 => x"822ea638",
   722 => x"71822689",
   723 => x"3871812e",
   724 => x"a93897cf",
   725 => x"0471832e",
   726 => x"b1387184",
   727 => x"2e098106",
   728 => x"80ed3888",
   729 => x"1308518f",
   730 => x"a72d97cf",
   731 => x"04b9f408",
   732 => x"51881308",
   733 => x"52712d97",
   734 => x"cf04810b",
   735 => x"8814082b",
   736 => x"b9e00832",
   737 => x"b9e00c97",
   738 => x"a5048813",
   739 => x"80f52d81",
   740 => x"058b1480",
   741 => x"f52d5354",
   742 => x"71742483",
   743 => x"38805473",
   744 => x"881481b7",
   745 => x"2d8e8c2d",
   746 => x"97cf0475",
   747 => x"08802ea2",
   748 => x"38750851",
   749 => x"8b8b2db9",
   750 => x"8c088106",
   751 => x"5271802e",
   752 => x"8b38b9f4",
   753 => x"08518416",
   754 => x"0852712d",
   755 => x"88165675",
   756 => x"da388054",
   757 => x"800bb9a0",
   758 => x"0c738f06",
   759 => x"b99c0ca0",
   760 => x"5273b9f4",
   761 => x"082e0981",
   762 => x"069838b9",
   763 => x"f008ff05",
   764 => x"74327009",
   765 => x"81057072",
   766 => x"079f2a91",
   767 => x"71315151",
   768 => x"53537151",
   769 => x"82f92d81",
   770 => x"14548e74",
   771 => x"25c638b7",
   772 => x"cc085271",
   773 => x"b98c0c02",
   774 => x"98050d04",
   775 => x"02f4050d",
   776 => x"d45281ff",
   777 => x"720c7108",
   778 => x"5381ff72",
   779 => x"0c72882b",
   780 => x"83fe8006",
   781 => x"72087081",
   782 => x"ff065152",
   783 => x"5381ff72",
   784 => x"0c727107",
   785 => x"882b7208",
   786 => x"7081ff06",
   787 => x"51525381",
   788 => x"ff720c72",
   789 => x"7107882b",
   790 => x"72087081",
   791 => x"ff067207",
   792 => x"b98c0c52",
   793 => x"53028c05",
   794 => x"0d0402f4",
   795 => x"050d7476",
   796 => x"7181ff06",
   797 => x"d40c5353",
   798 => x"b9fc0885",
   799 => x"3871892b",
   800 => x"5271982a",
   801 => x"d40c7190",
   802 => x"2a7081ff",
   803 => x"06d40c51",
   804 => x"71882a70",
   805 => x"81ff06d4",
   806 => x"0c517181",
   807 => x"ff06d40c",
   808 => x"72902a70",
   809 => x"81ff06d4",
   810 => x"0c51d408",
   811 => x"7081ff06",
   812 => x"515182b8",
   813 => x"bf527081",
   814 => x"ff2e0981",
   815 => x"06943881",
   816 => x"ff0bd40c",
   817 => x"d4087081",
   818 => x"ff06ff14",
   819 => x"54515171",
   820 => x"e53870b9",
   821 => x"8c0c028c",
   822 => x"050d0402",
   823 => x"fc050d81",
   824 => x"c75181ff",
   825 => x"0bd40cff",
   826 => x"11517080",
   827 => x"25f43802",
   828 => x"84050d04",
   829 => x"02f4050d",
   830 => x"81ff0bd4",
   831 => x"0c935380",
   832 => x"5287fc80",
   833 => x"c15198ea",
   834 => x"2db98c08",
   835 => x"8b3881ff",
   836 => x"0bd40c81",
   837 => x"539aa104",
   838 => x"99db2dff",
   839 => x"135372df",
   840 => x"3872b98c",
   841 => x"0c028c05",
   842 => x"0d0402ec",
   843 => x"050d810b",
   844 => x"b9fc0c84",
   845 => x"54d00870",
   846 => x"8f2a7081",
   847 => x"06515153",
   848 => x"72f33872",
   849 => x"d00c99db",
   850 => x"2db48851",
   851 => x"85fe2dd0",
   852 => x"08708f2a",
   853 => x"70810651",
   854 => x"515372f3",
   855 => x"38810bd0",
   856 => x"0cb15380",
   857 => x"5284d480",
   858 => x"c05198ea",
   859 => x"2db98c08",
   860 => x"812e9338",
   861 => x"72822ebd",
   862 => x"38ff1353",
   863 => x"72e538ff",
   864 => x"145473ff",
   865 => x"b03899db",
   866 => x"2d83aa52",
   867 => x"849c80c8",
   868 => x"5198ea2d",
   869 => x"b98c0881",
   870 => x"2e098106",
   871 => x"9238989c",
   872 => x"2db98c08",
   873 => x"83ffff06",
   874 => x"537283aa",
   875 => x"2e9d3899",
   876 => x"f42d9bc6",
   877 => x"04b49451",
   878 => x"85fe2d80",
   879 => x"539d9404",
   880 => x"b4ac5185",
   881 => x"fe2d8054",
   882 => x"9ce60481",
   883 => x"ff0bd40c",
   884 => x"b15499db",
   885 => x"2d8fcf53",
   886 => x"805287fc",
   887 => x"80f75198",
   888 => x"ea2db98c",
   889 => x"0855b98c",
   890 => x"08812e09",
   891 => x"81069b38",
   892 => x"81ff0bd4",
   893 => x"0c820a52",
   894 => x"849c80e9",
   895 => x"5198ea2d",
   896 => x"b98c0880",
   897 => x"2e8d3899",
   898 => x"db2dff13",
   899 => x"5372c938",
   900 => x"9cd90481",
   901 => x"ff0bd40c",
   902 => x"b98c0852",
   903 => x"87fc80fa",
   904 => x"5198ea2d",
   905 => x"b98c08b1",
   906 => x"3881ff0b",
   907 => x"d40cd408",
   908 => x"5381ff0b",
   909 => x"d40c81ff",
   910 => x"0bd40c81",
   911 => x"ff0bd40c",
   912 => x"81ff0bd4",
   913 => x"0c72862a",
   914 => x"70810676",
   915 => x"56515372",
   916 => x"9538b98c",
   917 => x"08549ce6",
   918 => x"0473822e",
   919 => x"fee238ff",
   920 => x"145473fe",
   921 => x"ed3873b9",
   922 => x"fc0c738b",
   923 => x"38815287",
   924 => x"fc80d051",
   925 => x"98ea2d81",
   926 => x"ff0bd40c",
   927 => x"d008708f",
   928 => x"2a708106",
   929 => x"51515372",
   930 => x"f33872d0",
   931 => x"0c81ff0b",
   932 => x"d40c8153",
   933 => x"72b98c0c",
   934 => x"0294050d",
   935 => x"0402e805",
   936 => x"0d785580",
   937 => x"5681ff0b",
   938 => x"d40cd008",
   939 => x"708f2a70",
   940 => x"81065151",
   941 => x"5372f338",
   942 => x"82810bd0",
   943 => x"0c81ff0b",
   944 => x"d40c7752",
   945 => x"87fc80d1",
   946 => x"5198ea2d",
   947 => x"80dbc6df",
   948 => x"54b98c08",
   949 => x"802e8a38",
   950 => x"b4cc5185",
   951 => x"fe2d9eb4",
   952 => x"0481ff0b",
   953 => x"d40cd408",
   954 => x"7081ff06",
   955 => x"51537281",
   956 => x"fe2e0981",
   957 => x"069d3880",
   958 => x"ff53989c",
   959 => x"2db98c08",
   960 => x"75708405",
   961 => x"570cff13",
   962 => x"53728025",
   963 => x"ed388156",
   964 => x"9e9904ff",
   965 => x"145473c9",
   966 => x"3881ff0b",
   967 => x"d40c81ff",
   968 => x"0bd40cd0",
   969 => x"08708f2a",
   970 => x"70810651",
   971 => x"515372f3",
   972 => x"3872d00c",
   973 => x"75b98c0c",
   974 => x"0298050d",
   975 => x"0402e805",
   976 => x"0d77797b",
   977 => x"58555580",
   978 => x"53727625",
   979 => x"a3387470",
   980 => x"81055680",
   981 => x"f52d7470",
   982 => x"81055680",
   983 => x"f52d5252",
   984 => x"71712e86",
   985 => x"3881519e",
   986 => x"f2048113",
   987 => x"539ec904",
   988 => x"805170b9",
   989 => x"8c0c0298",
   990 => x"050d0402",
   991 => x"ec050d76",
   992 => x"5574802e",
   993 => x"be389a15",
   994 => x"80e02d51",
   995 => x"acb52db9",
   996 => x"8c08b98c",
   997 => x"0880c0b0",
   998 => x"0cb98c08",
   999 => x"545480c0",
  1000 => x"8c08802e",
  1001 => x"99389415",
  1002 => x"80e02d51",
  1003 => x"acb52db9",
  1004 => x"8c08902b",
  1005 => x"83fff00a",
  1006 => x"06707507",
  1007 => x"51537280",
  1008 => x"c0b00c80",
  1009 => x"c0b00853",
  1010 => x"72802e9d",
  1011 => x"3880c084",
  1012 => x"08fe1471",
  1013 => x"2980c098",
  1014 => x"080580c0",
  1015 => x"b40c7084",
  1016 => x"2b80c090",
  1017 => x"0c54a097",
  1018 => x"0480c09c",
  1019 => x"0880c0b0",
  1020 => x"0c80c0a0",
  1021 => x"0880c0b4",
  1022 => x"0c80c08c",
  1023 => x"08802e8b",
  1024 => x"3880c084",
  1025 => x"08842b53",
  1026 => x"a0920480",
  1027 => x"c0a40884",
  1028 => x"2b537280",
  1029 => x"c0900c02",
  1030 => x"94050d04",
  1031 => x"02d8050d",
  1032 => x"800b80c0",
  1033 => x"8c0c8454",
  1034 => x"9aaa2db9",
  1035 => x"8c08802e",
  1036 => x"9538ba80",
  1037 => x"5280519d",
  1038 => x"9d2db98c",
  1039 => x"08802e86",
  1040 => x"38fe54a0",
  1041 => x"ce04ff14",
  1042 => x"54738024",
  1043 => x"db38738c",
  1044 => x"38b4dc51",
  1045 => x"85fe2d73",
  1046 => x"55a5f004",
  1047 => x"8056810b",
  1048 => x"80c0b80c",
  1049 => x"8853b4f0",
  1050 => x"52bab651",
  1051 => x"9ebd2db9",
  1052 => x"8c08762e",
  1053 => x"09810688",
  1054 => x"38b98c08",
  1055 => x"80c0b80c",
  1056 => x"8853b4fc",
  1057 => x"52bad251",
  1058 => x"9ebd2db9",
  1059 => x"8c088838",
  1060 => x"b98c0880",
  1061 => x"c0b80c80",
  1062 => x"c0b80880",
  1063 => x"2e80f638",
  1064 => x"bdc60b80",
  1065 => x"f52dbdc7",
  1066 => x"0b80f52d",
  1067 => x"71982b71",
  1068 => x"902b07bd",
  1069 => x"c80b80f5",
  1070 => x"2d70882b",
  1071 => x"7207bdc9",
  1072 => x"0b80f52d",
  1073 => x"7107bdfe",
  1074 => x"0b80f52d",
  1075 => x"bdff0b80",
  1076 => x"f52d7188",
  1077 => x"2b07535f",
  1078 => x"54525a56",
  1079 => x"57557381",
  1080 => x"abaa2e09",
  1081 => x"81068d38",
  1082 => x"7551ac85",
  1083 => x"2db98c08",
  1084 => x"56a28104",
  1085 => x"7382d4d5",
  1086 => x"2e8738b5",
  1087 => x"8851a2c3",
  1088 => x"04ba8052",
  1089 => x"75519d9d",
  1090 => x"2db98c08",
  1091 => x"55b98c08",
  1092 => x"802e83dc",
  1093 => x"388853b4",
  1094 => x"fc52bad2",
  1095 => x"519ebd2d",
  1096 => x"b98c088a",
  1097 => x"38810b80",
  1098 => x"c08c0ca2",
  1099 => x"c9048853",
  1100 => x"b4f052ba",
  1101 => x"b6519ebd",
  1102 => x"2db98c08",
  1103 => x"802e8a38",
  1104 => x"b59c5185",
  1105 => x"fe2da3a3",
  1106 => x"04bdfe0b",
  1107 => x"80f52d54",
  1108 => x"7380d52e",
  1109 => x"09810680",
  1110 => x"ca38bdff",
  1111 => x"0b80f52d",
  1112 => x"547381aa",
  1113 => x"2e098106",
  1114 => x"ba38800b",
  1115 => x"ba800b80",
  1116 => x"f52d5654",
  1117 => x"7481e92e",
  1118 => x"83388154",
  1119 => x"7481eb2e",
  1120 => x"8c388055",
  1121 => x"73752e09",
  1122 => x"810682e4",
  1123 => x"38ba8b0b",
  1124 => x"80f52d55",
  1125 => x"748d38ba",
  1126 => x"8c0b80f5",
  1127 => x"2d547382",
  1128 => x"2e863880",
  1129 => x"55a5f004",
  1130 => x"ba8d0b80",
  1131 => x"f52d7080",
  1132 => x"c0840cff",
  1133 => x"0580c088",
  1134 => x"0cba8e0b",
  1135 => x"80f52dba",
  1136 => x"8f0b80f5",
  1137 => x"2d587605",
  1138 => x"77828029",
  1139 => x"057080c0",
  1140 => x"940cba90",
  1141 => x"0b80f52d",
  1142 => x"7080c0a8",
  1143 => x"0c80c08c",
  1144 => x"08595758",
  1145 => x"76802e81",
  1146 => x"ac388853",
  1147 => x"b4fc52ba",
  1148 => x"d2519ebd",
  1149 => x"2db98c08",
  1150 => x"81f63880",
  1151 => x"c0840870",
  1152 => x"842b80c0",
  1153 => x"900c7080",
  1154 => x"c0a40cba",
  1155 => x"a50b80f5",
  1156 => x"2dbaa40b",
  1157 => x"80f52d71",
  1158 => x"82802905",
  1159 => x"baa60b80",
  1160 => x"f52d7084",
  1161 => x"80802912",
  1162 => x"baa70b80",
  1163 => x"f52d7081",
  1164 => x"800a2912",
  1165 => x"7080c0ac",
  1166 => x"0c80c0a8",
  1167 => x"08712980",
  1168 => x"c0940805",
  1169 => x"7080c098",
  1170 => x"0cbaad0b",
  1171 => x"80f52dba",
  1172 => x"ac0b80f5",
  1173 => x"2d718280",
  1174 => x"2905baae",
  1175 => x"0b80f52d",
  1176 => x"70848080",
  1177 => x"2912baaf",
  1178 => x"0b80f52d",
  1179 => x"70982b81",
  1180 => x"f00a0672",
  1181 => x"057080c0",
  1182 => x"9c0cfe11",
  1183 => x"7e297705",
  1184 => x"80c0a00c",
  1185 => x"52595243",
  1186 => x"545e5152",
  1187 => x"59525d57",
  1188 => x"5957a5e9",
  1189 => x"04ba920b",
  1190 => x"80f52dba",
  1191 => x"910b80f5",
  1192 => x"2d718280",
  1193 => x"29057080",
  1194 => x"c0900c70",
  1195 => x"a02983ff",
  1196 => x"0570892a",
  1197 => x"7080c0a4",
  1198 => x"0cba970b",
  1199 => x"80f52dba",
  1200 => x"960b80f5",
  1201 => x"2d718280",
  1202 => x"29057080",
  1203 => x"c0ac0c7b",
  1204 => x"71291e70",
  1205 => x"80c0a00c",
  1206 => x"7d80c09c",
  1207 => x"0c730580",
  1208 => x"c0980c55",
  1209 => x"5e515155",
  1210 => x"5580519e",
  1211 => x"fb2d8155",
  1212 => x"74b98c0c",
  1213 => x"02a8050d",
  1214 => x"0402ec05",
  1215 => x"0d767087",
  1216 => x"2c7180ff",
  1217 => x"06555654",
  1218 => x"80c08c08",
  1219 => x"8a387388",
  1220 => x"2c7481ff",
  1221 => x"065455ba",
  1222 => x"805280c0",
  1223 => x"94081551",
  1224 => x"9d9d2db9",
  1225 => x"8c0854b9",
  1226 => x"8c08802e",
  1227 => x"b43880c0",
  1228 => x"8c08802e",
  1229 => x"98387284",
  1230 => x"29ba8005",
  1231 => x"70085253",
  1232 => x"ac852db9",
  1233 => x"8c08f00a",
  1234 => x"0653a6df",
  1235 => x"047210ba",
  1236 => x"80057080",
  1237 => x"e02d5253",
  1238 => x"acb52db9",
  1239 => x"8c085372",
  1240 => x"5473b98c",
  1241 => x"0c029405",
  1242 => x"0d0402e0",
  1243 => x"050d7970",
  1244 => x"842c80c0",
  1245 => x"b4080571",
  1246 => x"8f065255",
  1247 => x"53728938",
  1248 => x"ba805273",
  1249 => x"519d9d2d",
  1250 => x"72a029ba",
  1251 => x"80055480",
  1252 => x"7480f52d",
  1253 => x"56537473",
  1254 => x"2e833881",
  1255 => x"537481e5",
  1256 => x"2e81ef38",
  1257 => x"81707406",
  1258 => x"54587280",
  1259 => x"2e81e338",
  1260 => x"8b1480f5",
  1261 => x"2d70832a",
  1262 => x"79065856",
  1263 => x"769838b7",
  1264 => x"d0085372",
  1265 => x"883872be",
  1266 => x"800b81b7",
  1267 => x"2d76b7d0",
  1268 => x"0c7353a9",
  1269 => x"9404758f",
  1270 => x"2e098106",
  1271 => x"81b43874",
  1272 => x"9f068d29",
  1273 => x"bdf31151",
  1274 => x"53811480",
  1275 => x"f52d7370",
  1276 => x"81055581",
  1277 => x"b72d8314",
  1278 => x"80f52d73",
  1279 => x"70810555",
  1280 => x"81b72d85",
  1281 => x"1480f52d",
  1282 => x"73708105",
  1283 => x"5581b72d",
  1284 => x"871480f5",
  1285 => x"2d737081",
  1286 => x"055581b7",
  1287 => x"2d891480",
  1288 => x"f52d7370",
  1289 => x"81055581",
  1290 => x"b72d8e14",
  1291 => x"80f52d73",
  1292 => x"70810555",
  1293 => x"81b72d90",
  1294 => x"1480f52d",
  1295 => x"73708105",
  1296 => x"5581b72d",
  1297 => x"921480f5",
  1298 => x"2d737081",
  1299 => x"055581b7",
  1300 => x"2d941480",
  1301 => x"f52d7370",
  1302 => x"81055581",
  1303 => x"b72d9614",
  1304 => x"80f52d73",
  1305 => x"70810555",
  1306 => x"81b72d98",
  1307 => x"1480f52d",
  1308 => x"73708105",
  1309 => x"5581b72d",
  1310 => x"9c1480f5",
  1311 => x"2d737081",
  1312 => x"055581b7",
  1313 => x"2d9e1480",
  1314 => x"f52d7381",
  1315 => x"b72d77b7",
  1316 => x"d00c8053",
  1317 => x"72b98c0c",
  1318 => x"02a0050d",
  1319 => x"0402cc05",
  1320 => x"0d7e605e",
  1321 => x"5a800b80",
  1322 => x"c0b00880",
  1323 => x"c0b40859",
  1324 => x"5c568058",
  1325 => x"80c09008",
  1326 => x"782e81b0",
  1327 => x"38778f06",
  1328 => x"a0175754",
  1329 => x"738f38ba",
  1330 => x"80527651",
  1331 => x"8117579d",
  1332 => x"9d2dba80",
  1333 => x"56807680",
  1334 => x"f52d5654",
  1335 => x"74742e83",
  1336 => x"38815474",
  1337 => x"81e52e80",
  1338 => x"f7388170",
  1339 => x"7506555c",
  1340 => x"73802e80",
  1341 => x"eb388b16",
  1342 => x"80f52d98",
  1343 => x"06597880",
  1344 => x"df388b53",
  1345 => x"7c527551",
  1346 => x"9ebd2db9",
  1347 => x"8c0880d0",
  1348 => x"389c1608",
  1349 => x"51ac852d",
  1350 => x"b98c0884",
  1351 => x"1b0c9a16",
  1352 => x"80e02d51",
  1353 => x"acb52db9",
  1354 => x"8c08b98c",
  1355 => x"08881c0c",
  1356 => x"b98c0855",
  1357 => x"5580c08c",
  1358 => x"08802e98",
  1359 => x"38941680",
  1360 => x"e02d51ac",
  1361 => x"b52db98c",
  1362 => x"08902b83",
  1363 => x"fff00a06",
  1364 => x"70165154",
  1365 => x"73881b0c",
  1366 => x"787a0c7b",
  1367 => x"54aba504",
  1368 => x"81185880",
  1369 => x"c0900878",
  1370 => x"26fed238",
  1371 => x"80c08c08",
  1372 => x"802eb038",
  1373 => x"7a51a5f9",
  1374 => x"2db98c08",
  1375 => x"b98c0880",
  1376 => x"fffffff8",
  1377 => x"06555b73",
  1378 => x"80ffffff",
  1379 => x"f82e9438",
  1380 => x"b98c08fe",
  1381 => x"0580c084",
  1382 => x"082980c0",
  1383 => x"98080557",
  1384 => x"a9b20480",
  1385 => x"5473b98c",
  1386 => x"0c02b405",
  1387 => x"0d0402f4",
  1388 => x"050d7470",
  1389 => x"08810571",
  1390 => x"0c700880",
  1391 => x"c0880806",
  1392 => x"5353718e",
  1393 => x"38881308",
  1394 => x"51a5f92d",
  1395 => x"b98c0888",
  1396 => x"140c810b",
  1397 => x"b98c0c02",
  1398 => x"8c050d04",
  1399 => x"02f0050d",
  1400 => x"75881108",
  1401 => x"fe0580c0",
  1402 => x"84082980",
  1403 => x"c0980811",
  1404 => x"720880c0",
  1405 => x"88080605",
  1406 => x"79555354",
  1407 => x"549d9d2d",
  1408 => x"0290050d",
  1409 => x"0402f405",
  1410 => x"0d747088",
  1411 => x"2a83fe80",
  1412 => x"06707298",
  1413 => x"2a077288",
  1414 => x"2b87fc80",
  1415 => x"80067398",
  1416 => x"2b81f00a",
  1417 => x"06717307",
  1418 => x"07b98c0c",
  1419 => x"56515351",
  1420 => x"028c050d",
  1421 => x"0402f805",
  1422 => x"0d028e05",
  1423 => x"80f52d74",
  1424 => x"882b0770",
  1425 => x"83ffff06",
  1426 => x"b98c0c51",
  1427 => x"0288050d",
  1428 => x"0402f405",
  1429 => x"0d747678",
  1430 => x"53545280",
  1431 => x"71259738",
  1432 => x"72708105",
  1433 => x"5480f52d",
  1434 => x"72708105",
  1435 => x"5481b72d",
  1436 => x"ff115170",
  1437 => x"eb388072",
  1438 => x"81b72d02",
  1439 => x"8c050d04",
  1440 => x"02e8050d",
  1441 => x"77568070",
  1442 => x"56547376",
  1443 => x"24b33880",
  1444 => x"c0900874",
  1445 => x"2eab3873",
  1446 => x"51a6ea2d",
  1447 => x"b98c08b9",
  1448 => x"8c080981",
  1449 => x"0570b98c",
  1450 => x"08079f2a",
  1451 => x"77058117",
  1452 => x"57575353",
  1453 => x"74762489",
  1454 => x"3880c090",
  1455 => x"087426d7",
  1456 => x"3872b98c",
  1457 => x"0c029805",
  1458 => x"0d0402f0",
  1459 => x"050db988",
  1460 => x"081651ad",
  1461 => x"802db98c",
  1462 => x"08802e9c",
  1463 => x"388b53b9",
  1464 => x"8c0852be",
  1465 => x"8051acd1",
  1466 => x"2d80c0bc",
  1467 => x"08547380",
  1468 => x"2e8638be",
  1469 => x"8051732d",
  1470 => x"0290050d",
  1471 => x"0402dc05",
  1472 => x"0d80705a",
  1473 => x"5574b988",
  1474 => x"0825b138",
  1475 => x"80c09008",
  1476 => x"752ea938",
  1477 => x"7851a6ea",
  1478 => x"2db98c08",
  1479 => x"09810570",
  1480 => x"b98c0807",
  1481 => x"9f2a7605",
  1482 => x"811b5b56",
  1483 => x"5474b988",
  1484 => x"08258938",
  1485 => x"80c09008",
  1486 => x"7926d938",
  1487 => x"80557880",
  1488 => x"c0900827",
  1489 => x"81d13878",
  1490 => x"51a6ea2d",
  1491 => x"b98c0880",
  1492 => x"2e81a538",
  1493 => x"b98c088b",
  1494 => x"0580f52d",
  1495 => x"70842a70",
  1496 => x"81067710",
  1497 => x"78842bbe",
  1498 => x"800b80f5",
  1499 => x"2d5c5c53",
  1500 => x"51555673",
  1501 => x"802e80c8",
  1502 => x"38741682",
  1503 => x"2bb0bb0b",
  1504 => x"b7dc120c",
  1505 => x"54777531",
  1506 => x"1080c0c0",
  1507 => x"11555690",
  1508 => x"74708105",
  1509 => x"5681b72d",
  1510 => x"a07481b7",
  1511 => x"2d7681ff",
  1512 => x"06811658",
  1513 => x"5473802e",
  1514 => x"89389c53",
  1515 => x"be8052af",
  1516 => x"b8048b53",
  1517 => x"b98c0852",
  1518 => x"80c0c216",
  1519 => x"51aff004",
  1520 => x"7416822b",
  1521 => x"adca0bb7",
  1522 => x"dc120c54",
  1523 => x"7681ff06",
  1524 => x"81165854",
  1525 => x"73802e89",
  1526 => x"389c53be",
  1527 => x"8052afe7",
  1528 => x"048b53b9",
  1529 => x"8c085277",
  1530 => x"75311080",
  1531 => x"c0c00551",
  1532 => x"7655acd1",
  1533 => x"2db08c04",
  1534 => x"74902975",
  1535 => x"31701080",
  1536 => x"c0c00551",
  1537 => x"54b98c08",
  1538 => x"7481b72d",
  1539 => x"81195974",
  1540 => x"8b24a338",
  1541 => x"aebe0474",
  1542 => x"90297531",
  1543 => x"701080c0",
  1544 => x"c0058c77",
  1545 => x"31575154",
  1546 => x"807481b7",
  1547 => x"2d9e14ff",
  1548 => x"16565474",
  1549 => x"f33802a4",
  1550 => x"050d0402",
  1551 => x"fc050db9",
  1552 => x"88081351",
  1553 => x"ad802db9",
  1554 => x"8c08802e",
  1555 => x"8838b98c",
  1556 => x"08519efb",
  1557 => x"2d800bb9",
  1558 => x"880cadfd",
  1559 => x"2d8e8c2d",
  1560 => x"0284050d",
  1561 => x"0402fc05",
  1562 => x"0d725170",
  1563 => x"fd2ead38",
  1564 => x"70fd248a",
  1565 => x"3870fc2e",
  1566 => x"80c438b1",
  1567 => x"c60470fe",
  1568 => x"2eb13870",
  1569 => x"ff2e0981",
  1570 => x"06bc38b9",
  1571 => x"88085170",
  1572 => x"802eb338",
  1573 => x"ff11b988",
  1574 => x"0cb1c604",
  1575 => x"b98808f0",
  1576 => x"0570b988",
  1577 => x"0c517080",
  1578 => x"259c3880",
  1579 => x"0bb9880c",
  1580 => x"b1c604b9",
  1581 => x"88088105",
  1582 => x"b9880cb1",
  1583 => x"c604b988",
  1584 => x"089005b9",
  1585 => x"880cadfd",
  1586 => x"2d8e8c2d",
  1587 => x"0284050d",
  1588 => x"0402fc05",
  1589 => x"0d800bb9",
  1590 => x"880cadfd",
  1591 => x"2d8d912d",
  1592 => x"b98c08b8",
  1593 => x"f80cb7d4",
  1594 => x"518fa72d",
  1595 => x"0284050d",
  1596 => x"047180c0",
  1597 => x"bc0c0400",
  1598 => x"00ffffff",
  1599 => x"ff00ffff",
  1600 => x"ffff00ff",
  1601 => x"ffffff00",
  1602 => x"52657365",
  1603 => x"74000000",
  1604 => x"52474220",
  1605 => x"5363616c",
  1606 => x"696e6720",
  1607 => x"10000000",
  1608 => x"5363616e",
  1609 => x"6c696e65",
  1610 => x"73000000",
  1611 => x"416e696d",
  1612 => x"61746500",
  1613 => x"4c6f6164",
  1614 => x"20696d61",
  1615 => x"67652010",
  1616 => x"00000000",
  1617 => x"45786974",
  1618 => x"00000000",
  1619 => x"54657374",
  1620 => x"20706174",
  1621 => x"7465726e",
  1622 => x"20310000",
  1623 => x"54657374",
  1624 => x"20706174",
  1625 => x"7465726e",
  1626 => x"20320000",
  1627 => x"54657374",
  1628 => x"20706174",
  1629 => x"7465726e",
  1630 => x"20330000",
  1631 => x"54657374",
  1632 => x"20706174",
  1633 => x"7465726e",
  1634 => x"20340000",
  1635 => x"52656400",
  1636 => x"47726565",
  1637 => x"6e000000",
  1638 => x"426c7565",
  1639 => x"00000000",
  1640 => x"496e6974",
  1641 => x"69616c20",
  1642 => x"524f4d20",
  1643 => x"6c6f6164",
  1644 => x"696e6720",
  1645 => x"6661696c",
  1646 => x"65640000",
  1647 => x"4f4b0000",
  1648 => x"496e6974",
  1649 => x"69616c69",
  1650 => x"7a696e67",
  1651 => x"20534420",
  1652 => x"63617264",
  1653 => x"0a000000",
  1654 => x"4c6f6164",
  1655 => x"696e6720",
  1656 => x"696e6974",
  1657 => x"69616c20",
  1658 => x"524f4d2e",
  1659 => x"2e2e0a00",
  1660 => x"50494331",
  1661 => x"20202020",
  1662 => x"52415700",
  1663 => x"16200000",
  1664 => x"14200000",
  1665 => x"15200000",
  1666 => x"53442069",
  1667 => x"6e69742e",
  1668 => x"2e2e0a00",
  1669 => x"53442063",
  1670 => x"61726420",
  1671 => x"72657365",
  1672 => x"74206661",
  1673 => x"696c6564",
  1674 => x"210a0000",
  1675 => x"53444843",
  1676 => x"20657272",
  1677 => x"6f72210a",
  1678 => x"00000000",
  1679 => x"57726974",
  1680 => x"65206661",
  1681 => x"696c6564",
  1682 => x"0a000000",
  1683 => x"52656164",
  1684 => x"20666169",
  1685 => x"6c65640a",
  1686 => x"00000000",
  1687 => x"43617264",
  1688 => x"20696e69",
  1689 => x"74206661",
  1690 => x"696c6564",
  1691 => x"0a000000",
  1692 => x"46415431",
  1693 => x"36202020",
  1694 => x"00000000",
  1695 => x"46415433",
  1696 => x"32202020",
  1697 => x"00000000",
  1698 => x"4e6f2070",
  1699 => x"61727469",
  1700 => x"74696f6e",
  1701 => x"20736967",
  1702 => x"0a000000",
  1703 => x"42616420",
  1704 => x"70617274",
  1705 => x"0a000000",
  1706 => x"4261636b",
  1707 => x"00000000",
  1708 => x"00000002",
  1709 => x"00000002",
  1710 => x"00001908",
  1711 => x"00000352",
  1712 => x"00000003",
  1713 => x"00001b14",
  1714 => x"00000004",
  1715 => x"00000004",
  1716 => x"00001910",
  1717 => x"00001b24",
  1718 => x"00000001",
  1719 => x"00001920",
  1720 => x"00000000",
  1721 => x"00000002",
  1722 => x"0000192c",
  1723 => x"00000324",
  1724 => x"00000002",
  1725 => x"00001934",
  1726 => x"000018d1",
  1727 => x"00000002",
  1728 => x"00001944",
  1729 => x"000006ab",
  1730 => x"00000000",
  1731 => x"00000000",
  1732 => x"00000000",
  1733 => x"0000194c",
  1734 => x"0000195c",
  1735 => x"0000196c",
  1736 => x"0000197c",
  1737 => x"00000005",
  1738 => x"0000198c",
  1739 => x"00000010",
  1740 => x"00000005",
  1741 => x"00001990",
  1742 => x"00000010",
  1743 => x"00000005",
  1744 => x"00001998",
  1745 => x"00000010",
  1746 => x"00000004",
  1747 => x"00001944",
  1748 => x"00001ab4",
  1749 => x"00000000",
  1750 => x"00000000",
  1751 => x"00000000",
  1752 => x"00000004",
  1753 => x"000019a0",
  1754 => x"00001b60",
  1755 => x"00000004",
  1756 => x"000019bc",
  1757 => x"00001ab4",
  1758 => x"00000000",
  1759 => x"00000000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000002",
  1782 => x"00002040",
  1783 => x"000016ca",
  1784 => x"00000002",
  1785 => x"0000205e",
  1786 => x"000016ca",
  1787 => x"00000002",
  1788 => x"0000207c",
  1789 => x"000016ca",
  1790 => x"00000002",
  1791 => x"0000209a",
  1792 => x"000016ca",
  1793 => x"00000002",
  1794 => x"000020b8",
  1795 => x"000016ca",
  1796 => x"00000002",
  1797 => x"000020d6",
  1798 => x"000016ca",
  1799 => x"00000002",
  1800 => x"000020f4",
  1801 => x"000016ca",
  1802 => x"00000002",
  1803 => x"00002112",
  1804 => x"000016ca",
  1805 => x"00000002",
  1806 => x"00002130",
  1807 => x"000016ca",
  1808 => x"00000002",
  1809 => x"0000214e",
  1810 => x"000016ca",
  1811 => x"00000002",
  1812 => x"0000216c",
  1813 => x"000016ca",
  1814 => x"00000002",
  1815 => x"0000218a",
  1816 => x"000016ca",
  1817 => x"00000002",
  1818 => x"000021a8",
  1819 => x"000016ca",
  1820 => x"00000004",
  1821 => x"00001aa8",
  1822 => x"00000000",
  1823 => x"00000000",
  1824 => x"00000000",
  1825 => x"00001865",
  1826 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

