-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0b98",
     9 => x"fc080b0b",
    10 => x"0b998008",
    11 => x"0b0b0b99",
    12 => x"84080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"99840c0b",
    16 => x"0b0b9980",
    17 => x"0c0b0b0b",
    18 => x"98fc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0b95e8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"98fc7099",
    57 => x"e0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"85fd0402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"998c0c9f",
    65 => x"0b99900c",
    66 => x"a0717081",
    67 => x"05533499",
    68 => x"9008ff05",
    69 => x"99900c99",
    70 => x"90088025",
    71 => x"eb38998c",
    72 => x"08ff0599",
    73 => x"8c0c998c",
    74 => x"088025d7",
    75 => x"38800b99",
    76 => x"900c800b",
    77 => x"998c0c02",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"998c0825",
    97 => x"8f3882bc",
    98 => x"2d998c08",
    99 => x"ff05998c",
   100 => x"0c82fe04",
   101 => x"998c0899",
   102 => x"90085351",
   103 => x"728a2e09",
   104 => x"8106b738",
   105 => x"7151719f",
   106 => x"24a03899",
   107 => x"8c08a029",
   108 => x"11f88011",
   109 => x"5151a071",
   110 => x"34999008",
   111 => x"81059990",
   112 => x"0c999008",
   113 => x"519f7125",
   114 => x"e238800b",
   115 => x"99900c99",
   116 => x"8c088105",
   117 => x"998c0c83",
   118 => x"ee0470a0",
   119 => x"2912f880",
   120 => x"11515172",
   121 => x"71349990",
   122 => x"08810599",
   123 => x"900c9990",
   124 => x"08a02e09",
   125 => x"81068e38",
   126 => x"800b9990",
   127 => x"0c998c08",
   128 => x"8105998c",
   129 => x"0c028c05",
   130 => x"0d0402ec",
   131 => x"050d800b",
   132 => x"99940cf6",
   133 => x"8c08f690",
   134 => x"0871882c",
   135 => x"565481ff",
   136 => x"06527372",
   137 => x"25883871",
   138 => x"54820b99",
   139 => x"940c7288",
   140 => x"2c7381ff",
   141 => x"06545574",
   142 => x"73258b38",
   143 => x"72999408",
   144 => x"84079994",
   145 => x"0c557384",
   146 => x"2b86a071",
   147 => x"25837131",
   148 => x"700b0b0b",
   149 => x"978c0c81",
   150 => x"712bff05",
   151 => x"f6880cfe",
   152 => x"cc13ff12",
   153 => x"2c788829",
   154 => x"ff940570",
   155 => x"812c9994",
   156 => x"08525852",
   157 => x"55515254",
   158 => x"76802e85",
   159 => x"38708107",
   160 => x"5170f694",
   161 => x"0c710981",
   162 => x"05f6800c",
   163 => x"72098105",
   164 => x"f6840c02",
   165 => x"94050d04",
   166 => x"02f4050d",
   167 => x"74537270",
   168 => x"81055480",
   169 => x"f52d5271",
   170 => x"802e8938",
   171 => x"715182f8",
   172 => x"2d859e04",
   173 => x"810b98fc",
   174 => x"0c028c05",
   175 => x"0d0402fc",
   176 => x"050d8af4",
   177 => x"2d80518a",
   178 => x"ae2d8aae",
   179 => x"2d8aae2d",
   180 => x"8aae2d70",
   181 => x"f00c70f4",
   182 => x"0c70f80c",
   183 => x"81115190",
   184 => x"7125e438",
   185 => x"8ae12d02",
   186 => x"84050d04",
   187 => x"02fc050d",
   188 => x"ec518371",
   189 => x"0c82710c",
   190 => x"0284050d",
   191 => x"0402f405",
   192 => x"0d810bec",
   193 => x"0c8ac92d",
   194 => x"87982d81",
   195 => x"f72d97cc",
   196 => x"518cf02d",
   197 => x"83528aae",
   198 => x"2d815184",
   199 => x"8a2dff12",
   200 => x"52718025",
   201 => x"f138880b",
   202 => x"97980b81",
   203 => x"b72d880b",
   204 => x"97a40b81",
   205 => x"b72d880b",
   206 => x"97b00b81",
   207 => x"b72d8ae1",
   208 => x"2d800bec",
   209 => x"0c87a42d",
   210 => x"8d802d97",
   211 => x"e00b80f5",
   212 => x"2d99c408",
   213 => x"81065353",
   214 => x"71802e85",
   215 => x"38728407",
   216 => x"5372fc0c",
   217 => x"97980b80",
   218 => x"f52df00c",
   219 => x"97a40b80",
   220 => x"f52df40c",
   221 => x"97b00b80",
   222 => x"f52df80c",
   223 => x"825298fc",
   224 => x"08853898",
   225 => x"fc085271",
   226 => x"ec0c86c5",
   227 => x"0471980c",
   228 => x"04ffb008",
   229 => x"98fc0c04",
   230 => x"810bffb0",
   231 => x"0c04800b",
   232 => x"ffb00c04",
   233 => x"02f4050d",
   234 => x"88a60498",
   235 => x"fc0881f0",
   236 => x"2e098106",
   237 => x"8938810b",
   238 => x"98f00c88",
   239 => x"a60498fc",
   240 => x"0881e02e",
   241 => x"09810689",
   242 => x"38810b98",
   243 => x"f40c88a6",
   244 => x"0498fc08",
   245 => x"5298f408",
   246 => x"802e8838",
   247 => x"98fc0881",
   248 => x"80055271",
   249 => x"842c728f",
   250 => x"06535398",
   251 => x"f008802e",
   252 => x"99387284",
   253 => x"2998b005",
   254 => x"72138171",
   255 => x"2b700973",
   256 => x"0806730c",
   257 => x"51535388",
   258 => x"9c047284",
   259 => x"2998b005",
   260 => x"72138371",
   261 => x"2b720807",
   262 => x"720c5353",
   263 => x"800b98f4",
   264 => x"0c800b98",
   265 => x"f00c9998",
   266 => x"5189a72d",
   267 => x"98fc08ff",
   268 => x"24fef838",
   269 => x"800b98fc",
   270 => x"0c028c05",
   271 => x"0d0402f8",
   272 => x"050d98b0",
   273 => x"528f5180",
   274 => x"72708405",
   275 => x"540cff11",
   276 => x"51708025",
   277 => x"f2380288",
   278 => x"050d0402",
   279 => x"f0050d75",
   280 => x"51879e2d",
   281 => x"70822cfc",
   282 => x"0698b011",
   283 => x"72109e06",
   284 => x"71087072",
   285 => x"2a708306",
   286 => x"82742b70",
   287 => x"09740676",
   288 => x"0c545156",
   289 => x"57535153",
   290 => x"87982d71",
   291 => x"98fc0c02",
   292 => x"90050d04",
   293 => x"02fc050d",
   294 => x"72518071",
   295 => x"0c800b84",
   296 => x"120c0284",
   297 => x"050d0402",
   298 => x"f0050d75",
   299 => x"70088412",
   300 => x"08535353",
   301 => x"ff547171",
   302 => x"2ea83887",
   303 => x"9e2d8413",
   304 => x"08708429",
   305 => x"14881170",
   306 => x"087081ff",
   307 => x"06841808",
   308 => x"81118706",
   309 => x"841a0c53",
   310 => x"51555151",
   311 => x"5187982d",
   312 => x"71547398",
   313 => x"fc0c0290",
   314 => x"050d0402",
   315 => x"f8050d87",
   316 => x"9e2de008",
   317 => x"708b2a70",
   318 => x"81065152",
   319 => x"5270802e",
   320 => x"9d389998",
   321 => x"08708429",
   322 => x"99a00573",
   323 => x"81ff0671",
   324 => x"0c515199",
   325 => x"98088111",
   326 => x"87069998",
   327 => x"0c51800b",
   328 => x"99c00c87",
   329 => x"912d8798",
   330 => x"2d028805",
   331 => x"0d0402fc",
   332 => x"050d879e",
   333 => x"2d810b99",
   334 => x"c00c8798",
   335 => x"2d99c008",
   336 => x"5170fa38",
   337 => x"0284050d",
   338 => x"0402fc05",
   339 => x"0d999851",
   340 => x"89942d88",
   341 => x"be2d89eb",
   342 => x"51878d2d",
   343 => x"0284050d",
   344 => x"0402fc05",
   345 => x"0d810b98",
   346 => x"f80c8151",
   347 => x"848a2d02",
   348 => x"84050d04",
   349 => x"02fc050d",
   350 => x"8afe0487",
   351 => x"a42d8751",
   352 => x"88db2d98",
   353 => x"fc08f438",
   354 => x"80da5188",
   355 => x"db2d98fc",
   356 => x"08e93898",
   357 => x"fc0898f8",
   358 => x"0c98fc08",
   359 => x"51848a2d",
   360 => x"0284050d",
   361 => x"0402ec05",
   362 => x"0d765480",
   363 => x"52870b88",
   364 => x"1580f52d",
   365 => x"56537472",
   366 => x"248338a0",
   367 => x"53725182",
   368 => x"f82d8112",
   369 => x"8b1580f5",
   370 => x"2d545272",
   371 => x"7225de38",
   372 => x"0294050d",
   373 => x"0402f005",
   374 => x"0d99d008",
   375 => x"5481f72d",
   376 => x"800b99d4",
   377 => x"0c730880",
   378 => x"2e818038",
   379 => x"820b9990",
   380 => x"0c99d408",
   381 => x"8f06998c",
   382 => x"0c730852",
   383 => x"71832e96",
   384 => x"38718326",
   385 => x"89387181",
   386 => x"2eaf388c",
   387 => x"d6047185",
   388 => x"2e9f388c",
   389 => x"d6048814",
   390 => x"80f52d84",
   391 => x"15089780",
   392 => x"53545285",
   393 => x"982d7184",
   394 => x"29137008",
   395 => x"52528cda",
   396 => x"0473518b",
   397 => x"a52d8cd6",
   398 => x"0499c408",
   399 => x"8815082c",
   400 => x"70810651",
   401 => x"5271802e",
   402 => x"87389784",
   403 => x"518cd304",
   404 => x"97885185",
   405 => x"982d8414",
   406 => x"08518598",
   407 => x"2d99d408",
   408 => x"810599d4",
   409 => x"0c8c1454",
   410 => x"8be50402",
   411 => x"90050d04",
   412 => x"7199d00c",
   413 => x"8bd52d99",
   414 => x"d408ff05",
   415 => x"99d80c04",
   416 => x"02e8050d",
   417 => x"99d00899",
   418 => x"dc085755",
   419 => x"875188db",
   420 => x"2d98fc08",
   421 => x"812a7081",
   422 => x"06515271",
   423 => x"802ea038",
   424 => x"8da60487",
   425 => x"a42d8751",
   426 => x"88db2d98",
   427 => x"fc08f438",
   428 => x"98f80881",
   429 => x"327098f8",
   430 => x"0c705252",
   431 => x"848a2d80",
   432 => x"0b99c80c",
   433 => x"800b99cc",
   434 => x"0c98f808",
   435 => x"82dd3880",
   436 => x"da5188db",
   437 => x"2d98fc08",
   438 => x"802e8a38",
   439 => x"99c80881",
   440 => x"800799c8",
   441 => x"0c80d951",
   442 => x"88db2d98",
   443 => x"fc08802e",
   444 => x"8a3899c8",
   445 => x"0880c007",
   446 => x"99c80c81",
   447 => x"945188db",
   448 => x"2d98fc08",
   449 => x"802e8938",
   450 => x"99c80890",
   451 => x"0799c80c",
   452 => x"81915188",
   453 => x"db2d98fc",
   454 => x"08802e89",
   455 => x"3899c808",
   456 => x"a00799c8",
   457 => x"0c81f551",
   458 => x"88db2d98",
   459 => x"fc08802e",
   460 => x"893899c8",
   461 => x"08810799",
   462 => x"c80c81f2",
   463 => x"5188db2d",
   464 => x"98fc0880",
   465 => x"2e893899",
   466 => x"c8088207",
   467 => x"99c80c81",
   468 => x"eb5188db",
   469 => x"2d98fc08",
   470 => x"802e8938",
   471 => x"99c80884",
   472 => x"0799c80c",
   473 => x"81f45188",
   474 => x"db2d98fc",
   475 => x"08802e89",
   476 => x"3899c808",
   477 => x"880799c8",
   478 => x"0c80d851",
   479 => x"88db2d98",
   480 => x"fc08802e",
   481 => x"8a3899cc",
   482 => x"08818007",
   483 => x"99cc0c92",
   484 => x"5188db2d",
   485 => x"98fc0880",
   486 => x"2e8a3899",
   487 => x"cc0880c0",
   488 => x"0799cc0c",
   489 => x"945188db",
   490 => x"2d98fc08",
   491 => x"802e8938",
   492 => x"99cc0890",
   493 => x"0799cc0c",
   494 => x"915188db",
   495 => x"2d98fc08",
   496 => x"802e8938",
   497 => x"99cc08a0",
   498 => x"0799cc0c",
   499 => x"9d5188db",
   500 => x"2d98fc08",
   501 => x"802e8938",
   502 => x"99cc0881",
   503 => x"0799cc0c",
   504 => x"9b5188db",
   505 => x"2d98fc08",
   506 => x"802e8938",
   507 => x"99cc0882",
   508 => x"0799cc0c",
   509 => x"9c5188db",
   510 => x"2d98fc08",
   511 => x"802e8938",
   512 => x"99cc0884",
   513 => x"0799cc0c",
   514 => x"a35188db",
   515 => x"2d98fc08",
   516 => x"802e8938",
   517 => x"99cc0888",
   518 => x"0799cc0c",
   519 => x"81fd5188",
   520 => x"db2d81fa",
   521 => x"5188db2d",
   522 => x"95dc0481",
   523 => x"f55188db",
   524 => x"2d98fc08",
   525 => x"812a7081",
   526 => x"06515271",
   527 => x"802eaf38",
   528 => x"99d80852",
   529 => x"71802e89",
   530 => x"38ff1299",
   531 => x"d80c90ee",
   532 => x"0499d408",
   533 => x"1099d408",
   534 => x"05708429",
   535 => x"16515288",
   536 => x"1208802e",
   537 => x"8938ff51",
   538 => x"88120852",
   539 => x"712d81f2",
   540 => x"5188db2d",
   541 => x"98fc0881",
   542 => x"2a708106",
   543 => x"51527180",
   544 => x"2eb13899",
   545 => x"d408ff11",
   546 => x"99d80856",
   547 => x"53537372",
   548 => x"25893881",
   549 => x"1499d80c",
   550 => x"91b30472",
   551 => x"10137084",
   552 => x"29165152",
   553 => x"88120880",
   554 => x"2e8938fe",
   555 => x"51881208",
   556 => x"52712d81",
   557 => x"fd5188db",
   558 => x"2d98fc08",
   559 => x"812a7081",
   560 => x"06515271",
   561 => x"802ead38",
   562 => x"99d80880",
   563 => x"2e893880",
   564 => x"0b99d80c",
   565 => x"91f40499",
   566 => x"d4081099",
   567 => x"d4080570",
   568 => x"84291651",
   569 => x"52881208",
   570 => x"802e8938",
   571 => x"fd518812",
   572 => x"0852712d",
   573 => x"81fa5188",
   574 => x"db2d98fc",
   575 => x"08812a70",
   576 => x"81065152",
   577 => x"71802eae",
   578 => x"3899d408",
   579 => x"ff115452",
   580 => x"99d80873",
   581 => x"25883872",
   582 => x"99d80c92",
   583 => x"b6047110",
   584 => x"12708429",
   585 => x"16515288",
   586 => x"1208802e",
   587 => x"8938fc51",
   588 => x"88120852",
   589 => x"712d99d8",
   590 => x"08705354",
   591 => x"73802e8a",
   592 => x"388c15ff",
   593 => x"15555592",
   594 => x"bc04820b",
   595 => x"99900c71",
   596 => x"8f06998c",
   597 => x"0c81eb51",
   598 => x"88db2d98",
   599 => x"fc08812a",
   600 => x"70810651",
   601 => x"5271802e",
   602 => x"ad387408",
   603 => x"852e0981",
   604 => x"06a43888",
   605 => x"1580f52d",
   606 => x"ff055271",
   607 => x"881681b7",
   608 => x"2d71982b",
   609 => x"52718025",
   610 => x"8838800b",
   611 => x"881681b7",
   612 => x"2d74518b",
   613 => x"a52d81f4",
   614 => x"5188db2d",
   615 => x"98fc0881",
   616 => x"2a708106",
   617 => x"51527180",
   618 => x"2eb33874",
   619 => x"08852e09",
   620 => x"8106aa38",
   621 => x"881580f5",
   622 => x"2d810552",
   623 => x"71881681",
   624 => x"b72d7181",
   625 => x"ff068b16",
   626 => x"80f52d54",
   627 => x"52727227",
   628 => x"87387288",
   629 => x"1681b72d",
   630 => x"74518ba5",
   631 => x"2d80da51",
   632 => x"88db2d98",
   633 => x"fc08812a",
   634 => x"70810651",
   635 => x"5271802e",
   636 => x"81a63899",
   637 => x"d00899d8",
   638 => x"08555373",
   639 => x"802e8a38",
   640 => x"8c13ff15",
   641 => x"555393fb",
   642 => x"04720852",
   643 => x"71822ea6",
   644 => x"38718226",
   645 => x"89387181",
   646 => x"2ea93895",
   647 => x"98047183",
   648 => x"2eb13871",
   649 => x"842e0981",
   650 => x"0680ed38",
   651 => x"88130851",
   652 => x"8cf02d95",
   653 => x"980499d8",
   654 => x"08518813",
   655 => x"0852712d",
   656 => x"95980481",
   657 => x"0b881408",
   658 => x"2b99c408",
   659 => x"3299c40c",
   660 => x"94ee0488",
   661 => x"1380f52d",
   662 => x"81058b14",
   663 => x"80f52d53",
   664 => x"54717424",
   665 => x"83388054",
   666 => x"73881481",
   667 => x"b72d8bd5",
   668 => x"2d959804",
   669 => x"7508802e",
   670 => x"a2387508",
   671 => x"5188db2d",
   672 => x"98fc0881",
   673 => x"06527180",
   674 => x"2e8b3899",
   675 => x"d8085184",
   676 => x"16085271",
   677 => x"2d881656",
   678 => x"75da3880",
   679 => x"54800b99",
   680 => x"900c738f",
   681 => x"06998c0c",
   682 => x"a0527399",
   683 => x"d8082e09",
   684 => x"81069838",
   685 => x"99d408ff",
   686 => x"05743270",
   687 => x"09810570",
   688 => x"72079f2a",
   689 => x"91713151",
   690 => x"51535371",
   691 => x"5182f82d",
   692 => x"8114548e",
   693 => x"7425c638",
   694 => x"98f80852",
   695 => x"7198fc0c",
   696 => x"0298050d",
   697 => x"04000000",
   698 => x"00ffffff",
   699 => x"ff00ffff",
   700 => x"ffff00ff",
   701 => x"ffffff00",
   702 => x"52656400",
   703 => x"47726565",
   704 => x"6e000000",
   705 => x"426c7565",
   706 => x"00000000",
   707 => x"45786974",
   708 => x"00000000",
   709 => x"52657365",
   710 => x"74000000",
   711 => x"52474220",
   712 => x"5363616c",
   713 => x"696e6720",
   714 => x"10000000",
   715 => x"5363616e",
   716 => x"6c696e65",
   717 => x"73000000",
   718 => x"416e696d",
   719 => x"61746500",
   720 => x"54657374",
   721 => x"20706174",
   722 => x"7465726e",
   723 => x"20310000",
   724 => x"54657374",
   725 => x"20706174",
   726 => x"7465726e",
   727 => x"20320000",
   728 => x"54657374",
   729 => x"20706174",
   730 => x"7465726e",
   731 => x"20330000",
   732 => x"54657374",
   733 => x"20706174",
   734 => x"7465726e",
   735 => x"20340000",
   736 => x"16200000",
   737 => x"14200000",
   738 => x"15200000",
   739 => x"00000002",
   740 => x"00000005",
   741 => x"00000af8",
   742 => x"00000010",
   743 => x"00000005",
   744 => x"00000afc",
   745 => x"00000010",
   746 => x"00000005",
   747 => x"00000b04",
   748 => x"00000010",
   749 => x"00000004",
   750 => x"00000b0c",
   751 => x"00000bcc",
   752 => x"00000000",
   753 => x"00000000",
   754 => x"00000000",
   755 => x"00000002",
   756 => x"00000b14",
   757 => x"000002ec",
   758 => x"00000003",
   759 => x"00000c20",
   760 => x"00000004",
   761 => x"00000004",
   762 => x"00000b1c",
   763 => x"00000b90",
   764 => x"00000001",
   765 => x"00000b2c",
   766 => x"00000000",
   767 => x"00000002",
   768 => x"00000b38",
   769 => x"000002be",
   770 => x"00000002",
   771 => x"00000b0c",
   772 => x"00000574",
   773 => x"00000000",
   774 => x"00000000",
   775 => x"00000000",
   776 => x"00000b40",
   777 => x"00000b50",
   778 => x"00000b60",
   779 => x"00000b70",
   780 => x"00000000",
   781 => x"00000000",
   782 => x"00000000",
   783 => x"00000000",
   784 => x"00000000",
   785 => x"00000000",
   786 => x"00000000",
   787 => x"00000000",
   788 => x"00000000",
   789 => x"00000000",
   790 => x"00000000",
   791 => x"00000000",
   792 => x"00000000",
   793 => x"00000000",
   794 => x"00000000",
   795 => x"00000000",
   796 => x"00000000",
   797 => x"00000000",
   798 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

